cfg[0] = { 1'b0, 8'h40, 8'h0}; // CH=0 OP=0
cfg[1] = { 1'b0, 8'h41, 8'h1}; // CH=1 OP=0
cfg[2] = { 1'b0, 8'h42, 8'h2}; // CH=2 OP=0
cfg[3] = { 1'b1, 8'h40, 8'h3}; // CH=3 OP=0
cfg[4] = { 1'b1, 8'h41, 8'h4}; // CH=4 OP=0
cfg[5] = { 1'b1, 8'h42, 8'h5}; // CH=5 OP=0
cfg[6] = { 1'b0, 8'h44, 8'h6}; // CH=0 OP=1
cfg[7] = { 1'b0, 8'h45, 8'h7}; // CH=1 OP=1
cfg[8] = { 1'b0, 8'h46, 8'h8}; // CH=2 OP=1
cfg[9] = { 1'b1, 8'h44, 8'h9}; // CH=3 OP=1
cfg[10] = { 1'b1, 8'h45, 8'ha}; // CH=4 OP=1
cfg[11] = { 1'b1, 8'h46, 8'hb}; // CH=5 OP=1
cfg[12] = { 1'b0, 8'h48, 8'hc}; // CH=0 OP=2
cfg[13] = { 1'b0, 8'h49, 8'hd}; // CH=1 OP=2
cfg[14] = { 1'b0, 8'h4a, 8'he}; // CH=2 OP=2
cfg[15] = { 1'b1, 8'h48, 8'hf}; // CH=3 OP=2
cfg[16] = { 1'b1, 8'h49, 8'h10}; // CH=4 OP=2
cfg[17] = { 1'b1, 8'h4a, 8'h11}; // CH=5 OP=2
cfg[18] = { 1'b0, 8'h4c, 8'h12}; // CH=0 OP=3
cfg[19] = { 1'b0, 8'h4d, 8'h13}; // CH=1 OP=3
cfg[20] = { 1'b0, 8'h4e, 8'h14}; // CH=2 OP=3
cfg[21] = { 1'b1, 8'h4c, 8'h15}; // CH=3 OP=3
cfg[22] = { 1'b1, 8'h4d, 8'h16}; // CH=4 OP=3
cfg[23] = { 1'b1, 8'h4e, 8'h17}; // CH=5 OP=3

cfg[24] = { 1'b0, 8'h0, 8'h00 }; // done
