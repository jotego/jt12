cfg[0] = { 1'b0, 8'h30, 8'h0}; // CH=0 OP=0
cfg[1] = { 1'b0, 8'h34, 8'h1}; // CH=0 OP=1
cfg[2] = { 1'b0, 8'h38, 8'h2}; // CH=0 OP=2
cfg[3] = { 1'b0, 8'h3c, 8'h3}; // CH=0 OP=3
cfg[4] = { 1'b0, 8'h31, 8'h4}; // CH=1 OP=0
cfg[5] = { 1'b0, 8'h35, 8'h5}; // CH=1 OP=1
cfg[6] = { 1'b0, 8'h39, 8'h6}; // CH=1 OP=2
cfg[7] = { 1'b0, 8'h3d, 8'h7}; // CH=1 OP=3
cfg[8] = { 1'b0, 8'h32, 8'h8}; // CH=2 OP=0
cfg[9] = { 1'b0, 8'h36, 8'h9}; // CH=2 OP=1
cfg[10] = { 1'b0, 8'h3a, 8'ha}; // CH=2 OP=2
cfg[11] = { 1'b0, 8'h3e, 8'hb}; // CH=2 OP=3
cfg[12] = { 1'b1, 8'h30, 8'hc}; // CH=3 OP=0
cfg[13] = { 1'b1, 8'h34, 8'hd}; // CH=3 OP=1
cfg[14] = { 1'b1, 8'h38, 8'he}; // CH=3 OP=2
cfg[15] = { 1'b1, 8'h3c, 8'hf}; // CH=3 OP=3
cfg[16] = { 1'b1, 8'h31, 8'h10}; // CH=4 OP=0
cfg[17] = { 1'b1, 8'h35, 8'h11}; // CH=4 OP=1
cfg[18] = { 1'b1, 8'h39, 8'h12}; // CH=4 OP=2
cfg[19] = { 1'b1, 8'h3d, 8'h13}; // CH=4 OP=3
cfg[20] = { 1'b1, 8'h32, 8'h14}; // CH=5 OP=0
cfg[21] = { 1'b1, 8'h36, 8'h15}; // CH=5 OP=1
cfg[22] = { 1'b1, 8'h3a, 8'h16}; // CH=5 OP=2
cfg[23] = { 1'b1, 8'h3e, 8'h17}; // CH=5 OP=3
cfg[24] = { 1'b0, 8'h40, 8'h18}; // CH=0 OP=0
cfg[25] = { 1'b0, 8'h44, 8'h19}; // CH=0 OP=1
cfg[26] = { 1'b0, 8'h48, 8'h1a}; // CH=0 OP=2
cfg[27] = { 1'b0, 8'h4c, 8'h1b}; // CH=0 OP=3
cfg[28] = { 1'b0, 8'h41, 8'h1c}; // CH=1 OP=0
cfg[29] = { 1'b0, 8'h45, 8'h1d}; // CH=1 OP=1
cfg[30] = { 1'b0, 8'h49, 8'h1e}; // CH=1 OP=2
cfg[31] = { 1'b0, 8'h4d, 8'h1f}; // CH=1 OP=3
cfg[32] = { 1'b0, 8'h42, 8'h20}; // CH=2 OP=0
cfg[33] = { 1'b0, 8'h46, 8'h21}; // CH=2 OP=1
cfg[34] = { 1'b0, 8'h4a, 8'h22}; // CH=2 OP=2
cfg[35] = { 1'b0, 8'h4e, 8'h23}; // CH=2 OP=3
cfg[36] = { 1'b1, 8'h40, 8'h24}; // CH=3 OP=0
cfg[37] = { 1'b1, 8'h44, 8'h25}; // CH=3 OP=1
cfg[38] = { 1'b1, 8'h48, 8'h26}; // CH=3 OP=2
cfg[39] = { 1'b1, 8'h4c, 8'h27}; // CH=3 OP=3
cfg[40] = { 1'b1, 8'h41, 8'h28}; // CH=4 OP=0
cfg[41] = { 1'b1, 8'h45, 8'h29}; // CH=4 OP=1
cfg[42] = { 1'b1, 8'h49, 8'h2a}; // CH=4 OP=2
cfg[43] = { 1'b1, 8'h4d, 8'h2b}; // CH=4 OP=3
cfg[44] = { 1'b1, 8'h42, 8'h2c}; // CH=5 OP=0
cfg[45] = { 1'b1, 8'h46, 8'h2d}; // CH=5 OP=1
cfg[46] = { 1'b1, 8'h4a, 8'h2e}; // CH=5 OP=2
cfg[47] = { 1'b1, 8'h4e, 8'h2f}; // CH=5 OP=3
cfg[48] = { 1'b0, 8'h50, 8'h30}; // CH=0 OP=0
cfg[49] = { 1'b0, 8'h54, 8'h31}; // CH=0 OP=1
cfg[50] = { 1'b0, 8'h58, 8'h32}; // CH=0 OP=2
cfg[51] = { 1'b0, 8'h5c, 8'h33}; // CH=0 OP=3
cfg[52] = { 1'b0, 8'h51, 8'h34}; // CH=1 OP=0
cfg[53] = { 1'b0, 8'h55, 8'h35}; // CH=1 OP=1
cfg[54] = { 1'b0, 8'h59, 8'h36}; // CH=1 OP=2
cfg[55] = { 1'b0, 8'h5d, 8'h37}; // CH=1 OP=3
cfg[56] = { 1'b0, 8'h52, 8'h38}; // CH=2 OP=0
cfg[57] = { 1'b0, 8'h56, 8'h39}; // CH=2 OP=1
cfg[58] = { 1'b0, 8'h5a, 8'h3a}; // CH=2 OP=2
cfg[59] = { 1'b0, 8'h5e, 8'h3b}; // CH=2 OP=3
cfg[60] = { 1'b1, 8'h50, 8'h3c}; // CH=3 OP=0
cfg[61] = { 1'b1, 8'h54, 8'h3d}; // CH=3 OP=1
cfg[62] = { 1'b1, 8'h58, 8'h3e}; // CH=3 OP=2
cfg[63] = { 1'b1, 8'h5c, 8'h3f}; // CH=3 OP=3
cfg[64] = { 1'b1, 8'h51, 8'h40}; // CH=4 OP=0
cfg[65] = { 1'b1, 8'h55, 8'h41}; // CH=4 OP=1
cfg[66] = { 1'b1, 8'h59, 8'h42}; // CH=4 OP=2
cfg[67] = { 1'b1, 8'h5d, 8'h43}; // CH=4 OP=3
cfg[68] = { 1'b1, 8'h52, 8'h44}; // CH=5 OP=0
cfg[69] = { 1'b1, 8'h56, 8'h45}; // CH=5 OP=1
cfg[70] = { 1'b1, 8'h5a, 8'h46}; // CH=5 OP=2
cfg[71] = { 1'b1, 8'h5e, 8'h47}; // CH=5 OP=3
cfg[72] = { 1'b0, 8'h60, 8'h48}; // CH=0 OP=0
cfg[73] = { 1'b0, 8'h64, 8'h49}; // CH=0 OP=1
cfg[74] = { 1'b0, 8'h68, 8'h4a}; // CH=0 OP=2
cfg[75] = { 1'b0, 8'h6c, 8'h4b}; // CH=0 OP=3
cfg[76] = { 1'b0, 8'h61, 8'h4c}; // CH=1 OP=0
cfg[77] = { 1'b0, 8'h65, 8'h4d}; // CH=1 OP=1
cfg[78] = { 1'b0, 8'h69, 8'h4e}; // CH=1 OP=2
cfg[79] = { 1'b0, 8'h6d, 8'h4f}; // CH=1 OP=3
cfg[80] = { 1'b0, 8'h62, 8'h50}; // CH=2 OP=0
cfg[81] = { 1'b0, 8'h66, 8'h51}; // CH=2 OP=1
cfg[82] = { 1'b0, 8'h6a, 8'h52}; // CH=2 OP=2
cfg[83] = { 1'b0, 8'h6e, 8'h53}; // CH=2 OP=3
cfg[84] = { 1'b1, 8'h60, 8'h54}; // CH=3 OP=0
cfg[85] = { 1'b1, 8'h64, 8'h55}; // CH=3 OP=1
cfg[86] = { 1'b1, 8'h68, 8'h56}; // CH=3 OP=2
cfg[87] = { 1'b1, 8'h6c, 8'h57}; // CH=3 OP=3
cfg[88] = { 1'b1, 8'h61, 8'h58}; // CH=4 OP=0
cfg[89] = { 1'b1, 8'h65, 8'h59}; // CH=4 OP=1
cfg[90] = { 1'b1, 8'h69, 8'h5a}; // CH=4 OP=2
cfg[91] = { 1'b1, 8'h6d, 8'h5b}; // CH=4 OP=3
cfg[92] = { 1'b1, 8'h62, 8'h5c}; // CH=5 OP=0
cfg[93] = { 1'b1, 8'h66, 8'h5d}; // CH=5 OP=1
cfg[94] = { 1'b1, 8'h6a, 8'h5e}; // CH=5 OP=2
cfg[95] = { 1'b1, 8'h6e, 8'h5f}; // CH=5 OP=3
cfg[96] = { 1'b0, 8'h70, 8'h60}; // CH=0 OP=0
cfg[97] = { 1'b0, 8'h74, 8'h61}; // CH=0 OP=1
cfg[98] = { 1'b0, 8'h78, 8'h62}; // CH=0 OP=2
cfg[99] = { 1'b0, 8'h7c, 8'h63}; // CH=0 OP=3
cfg[100] = { 1'b0, 8'h71, 8'h64}; // CH=1 OP=0
cfg[101] = { 1'b0, 8'h75, 8'h65}; // CH=1 OP=1
cfg[102] = { 1'b0, 8'h79, 8'h66}; // CH=1 OP=2
cfg[103] = { 1'b0, 8'h7d, 8'h67}; // CH=1 OP=3
cfg[104] = { 1'b0, 8'h72, 8'h68}; // CH=2 OP=0
cfg[105] = { 1'b0, 8'h76, 8'h69}; // CH=2 OP=1
cfg[106] = { 1'b0, 8'h7a, 8'h6a}; // CH=2 OP=2
cfg[107] = { 1'b0, 8'h7e, 8'h6b}; // CH=2 OP=3
cfg[108] = { 1'b1, 8'h70, 8'h6c}; // CH=3 OP=0
cfg[109] = { 1'b1, 8'h74, 8'h6d}; // CH=3 OP=1
cfg[110] = { 1'b1, 8'h78, 8'h6e}; // CH=3 OP=2
cfg[111] = { 1'b1, 8'h7c, 8'h6f}; // CH=3 OP=3
cfg[112] = { 1'b1, 8'h71, 8'h70}; // CH=4 OP=0
cfg[113] = { 1'b1, 8'h75, 8'h71}; // CH=4 OP=1
cfg[114] = { 1'b1, 8'h79, 8'h72}; // CH=4 OP=2
cfg[115] = { 1'b1, 8'h7d, 8'h73}; // CH=4 OP=3
cfg[116] = { 1'b1, 8'h72, 8'h74}; // CH=5 OP=0
cfg[117] = { 1'b1, 8'h76, 8'h75}; // CH=5 OP=1
cfg[118] = { 1'b1, 8'h7a, 8'h76}; // CH=5 OP=2
cfg[119] = { 1'b1, 8'h7e, 8'h77}; // CH=5 OP=3
cfg[120] = { 1'b0, 8'h80, 8'h78}; // CH=0 OP=0
cfg[121] = { 1'b0, 8'h84, 8'h79}; // CH=0 OP=1
cfg[122] = { 1'b0, 8'h88, 8'h7a}; // CH=0 OP=2
cfg[123] = { 1'b0, 8'h8c, 8'h7b}; // CH=0 OP=3
cfg[124] = { 1'b0, 8'h81, 8'h7c}; // CH=1 OP=0
cfg[125] = { 1'b0, 8'h85, 8'h7d}; // CH=1 OP=1
cfg[126] = { 1'b0, 8'h89, 8'h7e}; // CH=1 OP=2
cfg[127] = { 1'b0, 8'h8d, 8'h7f}; // CH=1 OP=3
cfg[128] = { 1'b0, 8'h82, 8'h80}; // CH=2 OP=0
cfg[129] = { 1'b0, 8'h86, 8'h81}; // CH=2 OP=1
cfg[130] = { 1'b0, 8'h8a, 8'h82}; // CH=2 OP=2
cfg[131] = { 1'b0, 8'h8e, 8'h83}; // CH=2 OP=3
cfg[132] = { 1'b1, 8'h80, 8'h84}; // CH=3 OP=0
cfg[133] = { 1'b1, 8'h84, 8'h85}; // CH=3 OP=1
cfg[134] = { 1'b1, 8'h88, 8'h86}; // CH=3 OP=2
cfg[135] = { 1'b1, 8'h8c, 8'h87}; // CH=3 OP=3
cfg[136] = { 1'b1, 8'h81, 8'h88}; // CH=4 OP=0
cfg[137] = { 1'b1, 8'h85, 8'h89}; // CH=4 OP=1
cfg[138] = { 1'b1, 8'h89, 8'h8a}; // CH=4 OP=2
cfg[139] = { 1'b1, 8'h8d, 8'h8b}; // CH=4 OP=3
cfg[140] = { 1'b1, 8'h82, 8'h8c}; // CH=5 OP=0
cfg[141] = { 1'b1, 8'h86, 8'h8d}; // CH=5 OP=1
cfg[142] = { 1'b1, 8'h8a, 8'h8e}; // CH=5 OP=2
cfg[143] = { 1'b1, 8'h8e, 8'h8f}; // CH=5 OP=3
cfg[144] = { 1'b0, 8'h90, 8'h90}; // CH=0 OP=0
cfg[145] = { 1'b0, 8'h94, 8'h91}; // CH=0 OP=1
cfg[146] = { 1'b0, 8'h98, 8'h92}; // CH=0 OP=2
cfg[147] = { 1'b0, 8'h9c, 8'h93}; // CH=0 OP=3
cfg[148] = { 1'b0, 8'h91, 8'h94}; // CH=1 OP=0
cfg[149] = { 1'b0, 8'h95, 8'h95}; // CH=1 OP=1
cfg[150] = { 1'b0, 8'h99, 8'h96}; // CH=1 OP=2
cfg[151] = { 1'b0, 8'h9d, 8'h97}; // CH=1 OP=3
cfg[152] = { 1'b0, 8'h92, 8'h98}; // CH=2 OP=0
cfg[153] = { 1'b0, 8'h96, 8'h99}; // CH=2 OP=1
cfg[154] = { 1'b0, 8'h9a, 8'h9a}; // CH=2 OP=2
cfg[155] = { 1'b0, 8'h9e, 8'h9b}; // CH=2 OP=3
cfg[156] = { 1'b1, 8'h90, 8'h9c}; // CH=3 OP=0
cfg[157] = { 1'b1, 8'h94, 8'h9d}; // CH=3 OP=1
cfg[158] = { 1'b1, 8'h98, 8'h9e}; // CH=3 OP=2
cfg[159] = { 1'b1, 8'h9c, 8'h9f}; // CH=3 OP=3
cfg[160] = { 1'b1, 8'h91, 8'ha0}; // CH=4 OP=0
cfg[161] = { 1'b1, 8'h95, 8'ha1}; // CH=4 OP=1
cfg[162] = { 1'b1, 8'h99, 8'ha2}; // CH=4 OP=2
cfg[163] = { 1'b1, 8'h9d, 8'ha3}; // CH=4 OP=3
cfg[164] = { 1'b1, 8'h92, 8'ha4}; // CH=5 OP=0
cfg[165] = { 1'b1, 8'h96, 8'ha5}; // CH=5 OP=1
cfg[166] = { 1'b1, 8'h9a, 8'ha6}; // CH=5 OP=2
cfg[167] = { 1'b1, 8'h9e, 8'ha7}; // CH=5 OP=3
cfg[168] = { 1'b0, 8'ha0, 8'ha8}; // CH=0 OP=0
cfg[169] = { 1'b0, 8'ha4, 8'ha9}; // CH=0 OP=1
cfg[170] = { 1'b0, 8'ha1, 8'haa}; // CH=1 OP=0
cfg[171] = { 1'b0, 8'ha5, 8'hab}; // CH=1 OP=1
cfg[172] = { 1'b0, 8'ha2, 8'hac}; // CH=2 OP=0
cfg[173] = { 1'b0, 8'ha6, 8'had}; // CH=2 OP=1
cfg[174] = { 1'b1, 8'ha0, 8'hae}; // CH=3 OP=0
cfg[175] = { 1'b1, 8'ha4, 8'haf}; // CH=3 OP=1
cfg[176] = { 1'b1, 8'ha1, 8'hb0}; // CH=4 OP=0
cfg[177] = { 1'b1, 8'ha5, 8'hb1}; // CH=4 OP=1
cfg[178] = { 1'b1, 8'ha2, 8'hb2}; // CH=5 OP=0
cfg[179] = { 1'b1, 8'ha6, 8'hb3}; // CH=5 OP=1
cfg[180] = { 1'b0, 8'hb0, 8'hb4}; // CH=0 OP=0
cfg[181] = { 1'b0, 8'hb4, 8'hb5}; // CH=0 OP=1
cfg[182] = { 1'b0, 8'hb1, 8'hb6}; // CH=1 OP=0
cfg[183] = { 1'b0, 8'hb5, 8'hb7}; // CH=1 OP=1
cfg[184] = { 1'b0, 8'hb2, 8'hb8}; // CH=2 OP=0
cfg[185] = { 1'b0, 8'hb6, 8'hb9}; // CH=2 OP=1
cfg[186] = { 1'b1, 8'hb0, 8'hba}; // CH=3 OP=0
cfg[187] = { 1'b1, 8'hb4, 8'hbb}; // CH=3 OP=1
cfg[188] = { 1'b1, 8'hb1, 8'hbc}; // CH=4 OP=0
cfg[189] = { 1'b1, 8'hb5, 8'hbd}; // CH=4 OP=1
cfg[190] = { 1'b1, 8'hb2, 8'hbe}; // CH=5 OP=0
cfg[191] = { 1'b1, 8'hb6, 8'hbf}; // CH=5 OP=1
cfg[192] = { 1'b0, 8'hc0, 8'hc0}; // CH=0 OP=0
cfg[193] = { 1'b0, 8'hc4, 8'hc1}; // CH=0 OP=1
cfg[194] = { 1'b0, 8'hc1, 8'hc2}; // CH=1 OP=0
cfg[195] = { 1'b0, 8'hc5, 8'hc3}; // CH=1 OP=1
cfg[196] = { 1'b0, 8'hc2, 8'hc4}; // CH=2 OP=0
cfg[197] = { 1'b0, 8'hc6, 8'hc5}; // CH=2 OP=1
cfg[198] = { 1'b1, 8'hc0, 8'hc6}; // CH=3 OP=0
cfg[199] = { 1'b1, 8'hc4, 8'hc7}; // CH=3 OP=1
cfg[200] = { 1'b1, 8'hc1, 8'hc8}; // CH=4 OP=0
cfg[201] = { 1'b1, 8'hc5, 8'hc9}; // CH=4 OP=1
cfg[202] = { 1'b1, 8'hc2, 8'hca}; // CH=5 OP=0
cfg[203] = { 1'b1, 8'hc6, 8'hcb}; // CH=5 OP=1

cfg[204] = { 1'b0, 8'h0, 8'h00 }; // done
