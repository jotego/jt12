cfg[0] = { 1'b1, 8'h69, 8'hc6}; // CH=4 OP=2
cfg[1] = { 1'b1, 8'hff, 8'h51}; // CH=6 OP=3
cfg[2] = { 1'b0, 8'hcd, 8'hec}; // CH=1 OP=3
cfg[3] = { 1'b0, 8'hf2, 8'hab}; // CH=2 OP=0
cfg[4] = { 1'b1, 8'h46, 8'he3}; // CH=5 OP=1
cfg[5] = { 1'b0, 8'h54, 8'hc2}; // CH=0 OP=1
cfg[6] = { 1'b0, 8'he8, 8'h1b}; // CH=0 OP=2
cfg[7] = { 1'b1, 8'h76, 8'h8d}; // CH=5 OP=1
cfg[8] = { 1'b0, 8'h63, 8'h2e}; // CH=3 OP=0
cfg[9] = { 1'b1, 8'hc9, 8'h9f}; // CH=4 OP=2
cfg[10] = { 1'b0, 8'h32, 8'h66}; // CH=2 OP=0
cfg[11] = { 1'b1, 8'h31, 8'hb7}; // CH=4 OP=0
cfg[12] = { 1'b0, 8'h5a, 8'ha3}; // CH=2 OP=2
cfg[13] = { 1'b1, 8'h58, 8'h5d}; // CH=3 OP=2
cfg[14] = { 1'b1, 8'hd4, 8'h5e}; // CH=3 OP=1
cfg[15] = { 1'b1, 8'hcd, 8'hb2}; // CH=4 OP=3
cfg[16] = { 1'b0, 8'hb4, 8'h9b}; // CH=0 OP=1
cfg[17] = { 1'b0, 8'h82, 8'h11}; // CH=2 OP=0
cfg[18] = { 1'b0, 8'h3d, 8'h41}; // CH=1 OP=3
cfg[19] = { 1'b0, 8'h70, 8'h87}; // CH=0 OP=0
cfg[20] = { 1'b1, 8'ha1, 8'h3e}; // CH=4 OP=0
cfg[21] = { 1'b1, 8'hfc, 8'he1}; // CH=3 OP=3
cfg[22] = { 1'b1, 8'h7e, 8'h3e}; // CH=5 OP=3
cfg[23] = { 1'b1, 8'hdc, 8'hea}; // CH=3 OP=3
cfg[24] = { 1'b1, 8'h8f, 8'h96}; // CH=6 OP=3
cfg[25] = { 1'b0, 8'hec, 8'h5c}; // CH=0 OP=3
cfg[26] = { 1'b0, 8'hfb, 8'h3b}; // CH=3 OP=2
cfg[27] = { 1'b0, 8'h3c, 8'haf}; // CH=0 OP=3
cfg[28] = { 1'b0, 8'hdb, 8'hec}; // CH=3 OP=2
cfg[29] = { 1'b0, 8'hfe, 8'h2}; // CH=2 OP=3
cfg[30] = { 1'b1, 8'hfa, 8'hfb}; // CH=5 OP=2
cfg[31] = { 1'b0, 8'hfb, 8'h3a}; // CH=3 OP=2
cfg[32] = { 1'b1, 8'he6, 8'hd1}; // CH=5 OP=1
cfg[33] = { 1'b1, 8'h7c, 8'h3c}; // CH=3 OP=3
cfg[34] = { 1'b0, 8'hd8, 8'h75}; // CH=0 OP=2
cfg[35] = { 1'b0, 8'h89, 8'h61}; // CH=1 OP=2
cfg[36] = { 1'b1, 8'hbb, 8'h5c}; // CH=6 OP=2
cfg[37] = { 1'b0, 8'h95, 8'h99}; // CH=1 OP=1
cfg[38] = { 1'b1, 8'hf1, 8'heb}; // CH=4 OP=0
cfg[39] = { 1'b1, 8'hef, 8'h5}; // CH=6 OP=3
cfg[40] = { 1'b1, 8'he9, 8'h0}; // CH=4 OP=2
cfg[41] = { 1'b1, 8'he5, 8'h3a}; // CH=4 OP=1
cfg[42] = { 1'b0, 8'hcb, 8'hb}; // CH=3 OP=2
cfg[43] = { 1'b0, 8'h47, 8'h48}; // CH=3 OP=1
cfg[44] = { 1'b0, 8'ha8, 8'hbd}; // CH=0 OP=2
cfg[45] = { 1'b0, 8'h64, 8'h7b}; // CH=0 OP=1
cfg[46] = { 1'b1, 8'h73, 8'h14}; // CH=6 OP=0
cfg[47] = { 1'b0, 8'h5e, 8'hc5}; // CH=2 OP=3
cfg[48] = { 1'b1, 8'h63, 8'h79}; // CH=6 OP=0
cfg[49] = { 1'b1, 8'h64, 8'h70}; // CH=3 OP=1
cfg[50] = { 1'b0, 8'h9e, 8'h11}; // CH=2 OP=3
cfg[51] = { 1'b1, 8'haa, 8'hdc}; // CH=5 OP=2
cfg[52] = { 1'b0, 8'hf2, 8'hac}; // CH=2 OP=0
cfg[53] = { 1'b1, 8'haf, 8'h10}; // CH=6 OP=3
cfg[54] = { 1'b1, 8'hcd, 8'h33}; // CH=4 OP=3
cfg[55] = { 1'b1, 8'h48, 8'h50}; // CH=3 OP=2
cfg[56] = { 1'b1, 8'h5c, 8'h15}; // CH=3 OP=3
cfg[57] = { 1'b1, 8'hba, 8'h6f}; // CH=5 OP=2
cfg[58] = { 1'b1, 8'hf5, 8'h7d}; // CH=4 OP=1
cfg[59] = { 1'b1, 8'h7f, 8'he1}; // CH=6 OP=3
cfg[60] = { 1'b1, 8'hf8, 8'hf8}; // CH=3 OP=2
cfg[61] = { 1'b0, 8'hb5, 8'h1b}; // CH=1 OP=1
cfg[62] = { 1'b0, 8'he8, 8'h4e}; // CH=0 OP=2
cfg[63] = { 1'b0, 8'h38, 8'h32}; // CH=0 OP=2
cfg[64] = { 1'b0, 8'h4d, 8'h79}; // CH=1 OP=3
cfg[65] = { 1'b1, 8'hbc, 8'h34}; // CH=3 OP=3
cfg[66] = { 1'b1, 8'h77, 8'h4e}; // CH=6 OP=1
cfg[67] = { 1'b0, 8'h6c, 8'hcb}; // CH=0 OP=3
cfg[68] = { 1'b1, 8'h86, 8'hac}; // CH=5 OP=1
cfg[69] = { 1'b1, 8'haa, 8'h2b}; // CH=5 OP=2
cfg[70] = { 1'b0, 8'ha2, 8'h55}; // CH=2 OP=0
cfg[71] = { 1'b0, 8'hb5, 8'h70}; // CH=1 OP=1
cfg[72] = { 1'b1, 8'h5c, 8'h3b}; // CH=3 OP=3
cfg[73] = { 1'b1, 8'h94, 8'h36}; // CH=3 OP=1
cfg[74] = { 1'b1, 8'he2, 8'haf}; // CH=5 OP=0
cfg[75] = { 1'b0, 8'h9e, 8'he4}; // CH=2 OP=3
cfg[76] = { 1'b1, 8'h49, 8'h32}; // CH=4 OP=2
cfg[77] = { 1'b1, 8'h4e, 8'h82}; // CH=5 OP=3
cfg[78] = { 1'b1, 8'h70, 8'h8}; // CH=3 OP=0
cfg[79] = { 1'b0, 8'h8a, 8'hb2}; // CH=2 OP=2
cfg[80] = { 1'b1, 8'h48, 8'h54}; // CH=3 OP=2
cfg[81] = { 1'b0, 8'hbc, 8'ha}; // CH=0 OP=3
cfg[82] = { 1'b1, 8'ha8, 8'he}; // CH=3 OP=2
cfg[83] = { 1'b0, 8'h5b, 8'hac}; // CH=3 OP=2
cfg[84] = { 1'b1, 8'h4c, 8'h8e}; // CH=3 OP=3
cfg[85] = { 1'b1, 8'h9b, 8'h2d}; // CH=6 OP=2
cfg[86] = { 1'b1, 8'he5, 8'h42}; // CH=4 OP=1
cfg[87] = { 1'b0, 8'h33, 8'hc4}; // CH=3 OP=0
cfg[88] = { 1'b1, 8'ha3, 8'hcd}; // CH=6 OP=0
cfg[89] = { 1'b0, 8'had, 8'h7f}; // CH=1 OP=3
cfg[90] = { 1'b0, 8'h47, 8'h76}; // CH=3 OP=1
cfg[91] = { 1'b0, 8'hec, 8'h32}; // CH=0 OP=3
cfg[92] = { 1'b0, 8'h30, 8'hc4}; // CH=0 OP=0
cfg[93] = { 1'b0, 8'h85, 8'h20}; // CH=1 OP=1
cfg[94] = { 1'b0, 8'hb2, 8'hfb}; // CH=2 OP=0
cfg[95] = { 1'b1, 8'hf4, 8'h4}; // CH=3 OP=1
cfg[96] = { 1'b0, 8'hb9, 8'hb}; // CH=1 OP=2
cfg[97] = { 1'b0, 8'h86, 8'hba}; // CH=2 OP=1
cfg[98] = { 1'b1, 8'hf1, 8'h3e}; // CH=4 OP=0
cfg[99] = { 1'b0, 8'h67, 8'hd9}; // CH=3 OP=1
cfg[100] = { 1'b1, 8'h99, 8'hb7}; // CH=4 OP=2
cfg[101] = { 1'b0, 8'he3, 8'ha3}; // CH=3 OP=0
cfg[102] = { 1'b0, 8'hd9, 8'hd3}; // CH=1 OP=2
cfg[103] = { 1'b0, 8'h5e, 8'hf7}; // CH=2 OP=3
cfg[104] = { 1'b0, 8'ha8, 8'hf2}; // CH=0 OP=2
cfg[105] = { 1'b0, 8'h94, 8'h5}; // CH=0 OP=1
cfg[106] = { 1'b1, 8'hb4, 8'hbe}; // CH=3 OP=1
cfg[107] = { 1'b0, 8'h78, 8'h44}; // CH=0 OP=2
cfg[108] = { 1'b0, 8'h69, 8'h49}; // CH=1 OP=2
cfg[109] = { 1'b0, 8'hd0, 8'h23}; // CH=0 OP=0
cfg[110] = { 1'b0, 8'h69, 8'hda}; // CH=1 OP=2
cfg[111] = { 1'b0, 8'h4c, 8'h7e}; // CH=0 OP=3
cfg[112] = { 1'b0, 8'hb3, 8'h51}; // CH=3 OP=0
cfg[113] = { 1'b0, 8'h53, 8'h84}; // CH=3 OP=0
cfg[114] = { 1'b0, 8'hfb, 8'h94}; // CH=3 OP=2
cfg[115] = { 1'b1, 8'h90, 8'h99}; // CH=3 OP=0
cfg[116] = { 1'b0, 8'h44, 8'h57}; // CH=0 OP=1
cfg[117] = { 1'b0, 8'hbc, 8'h9b}; // CH=0 OP=3
cfg[118] = { 1'b1, 8'hcf, 8'he5}; // CH=6 OP=3
cfg[119] = { 1'b0, 8'he9, 8'hf5}; // CH=1 OP=2
cfg[120] = { 1'b0, 8'h53, 8'h5e}; // CH=3 OP=0
cfg[121] = { 1'b0, 8'hd2, 8'haa}; // CH=2 OP=0
cfg[122] = { 1'b0, 8'h85, 8'hd0}; // CH=1 OP=1
cfg[123] = { 1'b0, 8'hd8, 8'h54}; // CH=0 OP=2
cfg[124] = { 1'b1, 8'hd4, 8'he8}; // CH=3 OP=1
cfg[125] = { 1'b0, 8'h64, 8'h82}; // CH=0 OP=1
cfg[126] = { 1'b0, 8'ha8, 8'hd9}; // CH=0 OP=2
cfg[127] = { 1'b1, 8'h65, 8'h75}; // CH=4 OP=1
cfg[128] = { 1'b0, 8'h8a, 8'h5a}; // CH=2 OP=2
cfg[129] = { 1'b1, 8'h80, 8'h62}; // CH=3 OP=0
cfg[130] = { 1'b1, 8'hde, 8'h44}; // CH=5 OP=3
cfg[131] = { 1'b0, 8'h89, 8'ha5}; // CH=1 OP=2
cfg[132] = { 1'b0, 8'h59, 8'h57}; // CH=1 OP=2
cfg[133] = { 1'b1, 8'had, 8'h51}; // CH=4 OP=3
cfg[134] = { 1'b0, 8'h95, 8'h86}; // CH=1 OP=1
cfg[135] = { 1'b0, 8'he4, 8'hec}; // CH=0 OP=1
cfg[136] = { 1'b1, 8'h8c, 8'hf1}; // CH=3 OP=3
cfg[137] = { 1'b0, 8'hf1, 8'h66}; // CH=1 OP=0
cfg[138] = { 1'b0, 8'h7c, 8'hc0}; // CH=0 OP=3
cfg[139] = { 1'b1, 8'hfc, 8'h22}; // CH=3 OP=3
cfg[140] = { 1'b0, 8'hda, 8'h66}; // CH=2 OP=2
cfg[141] = { 1'b1, 8'h63, 8'hb}; // CH=6 OP=0
cfg[142] = { 1'b1, 8'hbc, 8'h62}; // CH=3 OP=3
cfg[143] = { 1'b1, 8'h69, 8'hb4}; // CH=4 OP=2
cfg[144] = { 1'b1, 8'hff, 8'h3a}; // CH=6 OP=3
cfg[145] = { 1'b1, 8'h93, 8'h27}; // CH=6 OP=0
cfg[146] = { 1'b0, 8'hb8, 8'h7}; // CH=0 OP=2
cfg[147] = { 1'b1, 8'h34, 8'h11}; // CH=3 OP=1
cfg[148] = { 1'b1, 8'hef, 8'h8d}; // CH=6 OP=3
cfg[149] = { 1'b1, 8'hd4, 8'h89}; // CH=3 OP=1
cfg[150] = { 1'b0, 8'h35, 8'h63}; // CH=1 OP=1
cfg[151] = { 1'b1, 8'he4, 8'hc7}; // CH=3 OP=1
cfg[152] = { 1'b0, 8'h67, 8'h83}; // CH=3 OP=1
cfg[153] = { 1'b0, 8'h96, 8'hed}; // CH=2 OP=1
cfg[154] = { 1'b0, 8'h45, 8'hec}; // CH=1 OP=1
cfg[155] = { 1'b1, 8'hd8, 8'h2}; // CH=3 OP=2
cfg[156] = { 1'b1, 8'hf8, 8'ha}; // CH=3 OP=2
cfg[157] = { 1'b1, 8'hd1, 8'h77}; // CH=4 OP=0
cfg[158] = { 1'b1, 8'hc1, 8'h96}; // CH=4 OP=0
cfg[159] = { 1'b0, 8'h95, 8'h1f}; // CH=1 OP=1
cfg[160] = { 1'b0, 8'hca, 8'h82}; // CH=2 OP=2
cfg[161] = { 1'b0, 8'hae, 8'h49}; // CH=2 OP=3
cfg[162] = { 1'b0, 8'h68, 8'hcd}; // CH=0 OP=2
cfg[163] = { 1'b0, 8'h7a, 8'hac}; // CH=2 OP=2
cfg[164] = { 1'b0, 8'hb4, 8'hf2}; // CH=0 OP=1
cfg[165] = { 1'b0, 8'h99, 8'hca}; // CH=1 OP=2
cfg[166] = { 1'b0, 8'h37, 8'hc2}; // CH=3 OP=1
cfg[167] = { 1'b0, 8'hcf, 8'hcb}; // CH=3 OP=3
cfg[168] = { 1'b1, 8'hc3, 8'hc9}; // CH=6 OP=0
cfg[169] = { 1'b0, 8'h6e, 8'h5e}; // CH=2 OP=3
cfg[170] = { 1'b1, 8'hda, 8'h28}; // CH=5 OP=2
cfg[171] = { 1'b0, 8'h6a, 8'hd7}; // CH=2 OP=2
cfg[172] = { 1'b1, 8'hd2, 8'hed}; // CH=5 OP=0
cfg[173] = { 1'b1, 8'h4c, 8'h99}; // CH=3 OP=3
cfg[174] = { 1'b1, 8'h56, 8'h8b}; // CH=5 OP=1
cfg[175] = { 1'b0, 8'hd1, 8'hd4}; // CH=1 OP=0
cfg[176] = { 1'b0, 8'hd9, 8'he4}; // CH=1 OP=2
cfg[177] = { 1'b1, 8'ha3, 8'h45}; // CH=6 OP=0
cfg[178] = { 1'b1, 8'hff, 8'hc6}; // CH=6 OP=3
cfg[179] = { 1'b1, 8'hd9, 8'h2a}; // CH=4 OP=2
cfg[180] = { 1'b1, 8'h43, 8'h1}; // CH=6 OP=0
cfg[181] = { 1'b1, 8'h87, 8'hee}; // CH=6 OP=1
cfg[182] = { 1'b1, 8'h62, 8'h7c}; // CH=5 OP=0
cfg[183] = { 1'b0, 8'hfc, 8'h69}; // CH=0 OP=3
cfg[184] = { 1'b0, 8'hcd, 8'h81}; // CH=1 OP=3
cfg[185] = { 1'b1, 8'ha6, 8'h65}; // CH=5 OP=1
cfg[186] = { 1'b0, 8'h49, 8'hab}; // CH=1 OP=2
cfg[187] = { 1'b1, 8'h4b, 8'h71}; // CH=6 OP=2
cfg[188] = { 1'b0, 8'h75, 8'h3a}; // CH=1 OP=1
cfg[189] = { 1'b1, 8'h76, 8'h4f}; // CH=5 OP=1
cfg[190] = { 1'b0, 8'h64, 8'h7e}; // CH=0 OP=1
cfg[191] = { 1'b1, 8'heb, 8'h81}; // CH=6 OP=2
cfg[192] = { 1'b1, 8'hfe, 8'hfd}; // CH=5 OP=3
cfg[193] = { 1'b1, 8'h67, 8'h9b}; // CH=6 OP=1
cfg[194] = { 1'b1, 8'he9, 8'hd}; // CH=4 OP=2
cfg[195] = { 1'b0, 8'h4e, 8'h7e}; // CH=2 OP=3
cfg[196] = { 1'b0, 8'hf9, 8'hbd}; // CH=1 OP=2
cfg[197] = { 1'b0, 8'h6a, 8'h8c}; // CH=2 OP=2
cfg[198] = { 1'b1, 8'ha4, 8'h5b}; // CH=3 OP=1
cfg[199] = { 1'b0, 8'hf4, 8'h2}; // CH=0 OP=1
cfg[200] = { 1'b0, 8'h72, 8'hed}; // CH=2 OP=0
cfg[201] = { 1'b0, 8'hf3, 8'hec}; // CH=3 OP=0
cfg[202] = { 1'b1, 8'hf0, 8'h4d}; // CH=3 OP=0
cfg[203] = { 1'b0, 8'h8b, 8'h10}; // CH=3 OP=2
cfg[204] = { 1'b1, 8'h99, 8'hcf}; // CH=4 OP=2
cfg[205] = { 1'b0, 8'h9f, 8'h5b}; // CH=3 OP=3
cfg[206] = { 1'b0, 8'h98, 8'hd4}; // CH=0 OP=2
cfg[207] = { 1'b0, 8'hd1, 8'h61}; // CH=1 OP=0
cfg[208] = { 1'b0, 8'hbe, 8'ha7}; // CH=2 OP=3
cfg[209] = { 1'b1, 8'hab, 8'hbf}; // CH=6 OP=2
cfg[210] = { 1'b0, 8'h98, 8'hd5}; // CH=0 OP=2
cfg[211] = { 1'b1, 8'he5, 8'hd6}; // CH=4 OP=1
cfg[212] = { 1'b0, 8'hf6, 8'hd6}; // CH=2 OP=1
cfg[213] = { 1'b1, 8'hc5, 8'h3e}; // CH=4 OP=1
cfg[214] = { 1'b0, 8'haf, 8'h8e}; // CH=3 OP=3
cfg[215] = { 1'b0, 8'hb9, 8'hc6}; // CH=1 OP=2
cfg[216] = { 1'b1, 8'h8a, 8'hc9}; // CH=5 OP=2
cfg[217] = { 1'b1, 8'h97, 8'h70}; // CH=6 OP=1
cfg[218] = { 1'b0, 8'h56, 8'hc}; // CH=2 OP=1
cfg[219] = { 1'b1, 8'hd8, 8'h1a}; // CH=3 OP=2
cfg[220] = { 1'b1, 8'hc2, 8'h8b}; // CH=5 OP=0
cfg[221] = { 1'b1, 8'he3, 8'ha4}; // CH=6 OP=0
cfg[222] = { 1'b1, 8'h92, 8'hd2}; // CH=5 OP=0
cfg[223] = { 1'b0, 8'h4b, 8'h98}; // CH=3 OP=2
cfg[224] = { 1'b1, 8'hd5, 8'h61}; // CH=4 OP=1
cfg[225] = { 1'b1, 8'h6c, 8'hd1}; // CH=3 OP=3
cfg[226] = { 1'b1, 8'hc2, 8'hdd}; // CH=5 OP=0
cfg[227] = { 1'b0, 8'hed, 8'hf7}; // CH=1 OP=3
cfg[228] = { 1'b0, 8'hef, 8'h13}; // CH=3 OP=3
cfg[229] = { 1'b1, 8'hc7, 8'h20}; // CH=6 OP=1
cfg[230] = { 1'b0, 8'hdd, 8'hab}; // CH=1 OP=3
cfg[231] = { 1'b0, 8'h81, 8'h4d}; // CH=1 OP=0
cfg[232] = { 1'b0, 8'h53, 8'h1c}; // CH=3 OP=0
cfg[233] = { 1'b0, 8'heb, 8'hee}; // CH=3 OP=2
cfg[234] = { 1'b0, 8'h4c, 8'h24}; // CH=0 OP=3
cfg[235] = { 1'b1, 8'ha8, 8'h79}; // CH=3 OP=2
cfg[236] = { 1'b0, 8'h6a, 8'hfb}; // CH=2 OP=2
cfg[237] = { 1'b0, 8'h58, 8'hf3}; // CH=0 OP=2
cfg[238] = { 1'b0, 8'h47, 8'h6}; // CH=3 OP=1
cfg[239] = { 1'b1, 8'hd2, 8'h26}; // CH=5 OP=0
cfg[240] = { 1'b1, 8'h6c, 8'hb2}; // CH=3 OP=3
cfg[241] = { 1'b0, 8'hc0, 8'h3b}; // CH=0 OP=0
cfg[242] = { 1'b0, 8'hab, 8'h2a}; // CH=3 OP=2
cfg[243] = { 1'b0, 8'hf8, 8'h4e}; // CH=0 OP=2
cfg[244] = { 1'b0, 8'h9e, 8'hc7}; // CH=2 OP=3
cfg[245] = { 1'b1, 8'hdb, 8'h11}; // CH=6 OP=2
cfg[246] = { 1'b0, 8'ha7, 8'h60}; // CH=3 OP=1
cfg[247] = { 1'b1, 8'hb5, 8'h31}; // CH=4 OP=1
cfg[248] = { 1'b1, 8'ha0, 8'h3}; // CH=3 OP=0
cfg[249] = { 1'b1, 8'h47, 8'h22}; // CH=6 OP=1
cfg[250] = { 1'b1, 8'h9b, 8'hcd}; // CH=6 OP=2
cfg[251] = { 1'b1, 8'h56, 8'h78}; // CH=5 OP=1
cfg[252] = { 1'b1, 8'h4c, 8'h70}; // CH=3 OP=3
cfg[253] = { 1'b0, 8'hea, 8'h86}; // CH=2 OP=2
cfg[254] = { 1'b1, 8'hf2, 8'h98}; // CH=5 OP=0
cfg[255] = { 1'b1, 8'h53, 8'h9c}; // CH=6 OP=0
cfg[256] = { 1'b1, 8'hfa, 8'ha7}; // CH=5 OP=2
cfg[257] = { 1'b0, 8'hb0, 8'hd8}; // CH=0 OP=0
cfg[258] = { 1'b1, 8'h50, 8'hdb}; // CH=3 OP=0
cfg[259] = { 1'b0, 8'h5d, 8'hfd}; // CH=1 OP=3
cfg[260] = { 1'b1, 8'ha5, 8'h5a}; // CH=4 OP=1
cfg[261] = { 1'b0, 8'hfb, 8'ha3}; // CH=3 OP=2
cfg[262] = { 1'b1, 8'h47, 8'h13}; // CH=6 OP=1
cfg[263] = { 1'b0, 8'h31, 8'h9a}; // CH=1 OP=0
cfg[264] = { 1'b1, 8'h4e, 8'h32}; // CH=5 OP=3
cfg[265] = { 1'b0, 8'h5b, 8'h76}; // CH=3 OP=2
cfg[266] = { 1'b1, 8'hb6, 8'h71}; // CH=5 OP=1
cfg[267] = { 1'b1, 8'h6b, 8'h21}; // CH=6 OP=2
cfg[268] = { 1'b0, 8'hcf, 8'h71}; // CH=3 OP=3
cfg[269] = { 1'b1, 8'hf9, 8'h80}; // CH=4 OP=2
cfg[270] = { 1'b0, 8'h9c, 8'h62}; // CH=0 OP=3
cfg[271] = { 1'b1, 8'hb0, 8'h19}; // CH=3 OP=0
cfg[272] = { 1'b0, 8'h4a, 8'h6d}; // CH=2 OP=2
cfg[273] = { 1'b1, 8'h7c, 8'hd1}; // CH=3 OP=3
cfg[274] = { 1'b1, 8'h4a, 8'h1f}; // CH=5 OP=2
cfg[275] = { 1'b1, 8'hc0, 8'h7b}; // CH=3 OP=0
cfg[276] = { 1'b0, 8'h7b, 8'h31}; // CH=3 OP=2
cfg[277] = { 1'b0, 8'hed, 8'h36}; // CH=1 OP=3
cfg[278] = { 1'b0, 8'hbc, 8'h5b}; // CH=0 OP=3
cfg[279] = { 1'b0, 8'hb5, 8'hdb}; // CH=1 OP=1
cfg[280] = { 1'b0, 8'h52, 8'h3d}; // CH=2 OP=0
cfg[281] = { 1'b0, 8'hd4, 8'h57}; // CH=0 OP=1
cfg[282] = { 1'b0, 8'h95, 8'h4c}; // CH=1 OP=1
cfg[283] = { 1'b0, 8'hb5, 8'h97}; // CH=1 OP=1
cfg[284] = { 1'b0, 8'h30, 8'h80}; // CH=0 OP=0
cfg[285] = { 1'b0, 8'h61, 8'hdb}; // CH=1 OP=0
cfg[286] = { 1'b0, 8'hfd, 8'h56}; // CH=1 OP=3
cfg[287] = { 1'b0, 8'hc8, 8'h43}; // CH=0 OP=2
cfg[288] = { 1'b1, 8'hca, 8'hff}; // CH=5 OP=2
cfg[289] = { 1'b1, 8'ha8, 8'hb5}; // CH=3 OP=2
cfg[290] = { 1'b0, 8'h5e, 8'h7}; // CH=2 OP=3
cfg[291] = { 1'b1, 8'h33, 8'h9}; // CH=6 OP=0
cfg[292] = { 1'b0, 8'h57, 8'h55}; // CH=3 OP=1
cfg[293] = { 1'b1, 8'hee, 8'h1d}; // CH=5 OP=3
cfg[294] = { 1'b0, 8'h6e, 8'h2f}; // CH=2 OP=3
cfg[295] = { 1'b0, 8'h49, 8'h2}; // CH=1 OP=2
cfg[296] = { 1'b1, 8'ha0, 8'he2}; // CH=3 OP=0
cfg[297] = { 1'b1, 8'he3, 8'hf8}; // CH=6 OP=0
cfg[298] = { 1'b1, 8'he3, 8'h69}; // CH=6 OP=0
cfg[299] = { 1'b1, 8'h98, 8'hb6}; // CH=3 OP=2
cfg[300] = { 1'b1, 8'h9f, 8'h41}; // CH=6 OP=3
cfg[301] = { 1'b0, 8'ha8, 8'h22}; // CH=0 OP=2
cfg[302] = { 1'b1, 8'hfd, 8'hc8}; // CH=4 OP=3
cfg[303] = { 1'b0, 8'h90, 8'h4}; // CH=0 OP=0
cfg[304] = { 1'b0, 8'hfe, 8'h49}; // CH=2 OP=3
cfg[305] = { 1'b1, 8'h48, 8'h4b}; // CH=3 OP=2
cfg[306] = { 1'b0, 8'he8, 8'h2d}; // CH=0 OP=2
cfg[307] = { 1'b1, 8'hcb, 8'h25}; // CH=6 OP=2
cfg[308] = { 1'b0, 8'hae, 8'h8f}; // CH=2 OP=3
cfg[309] = { 1'b1, 8'h46, 8'h45}; // CH=5 OP=1
cfg[310] = { 1'b1, 8'he5, 8'h86}; // CH=4 OP=1
cfg[311] = { 1'b1, 8'h8d, 8'ha9}; // CH=4 OP=3
cfg[312] = { 1'b0, 8'h8a, 8'h71}; // CH=2 OP=2
cfg[313] = { 1'b0, 8'ha4, 8'h75}; // CH=0 OP=1
cfg[314] = { 1'b0, 8'hee, 8'h6a}; // CH=2 OP=3
cfg[315] = { 1'b0, 8'h39, 8'h7f}; // CH=1 OP=2
cfg[316] = { 1'b0, 8'h67, 8'h15}; // CH=3 OP=1
cfg[317] = { 1'b0, 8'h8c, 8'h2b}; // CH=0 OP=3
cfg[318] = { 1'b0, 8'h64, 8'h87}; // CH=0 OP=1
cfg[319] = { 1'b1, 8'hab, 8'h61}; // CH=6 OP=2
cfg[320] = { 1'b0, 8'h90, 8'he7}; // CH=0 OP=0
cfg[321] = { 1'b1, 8'he5, 8'h90}; // CH=4 OP=1
cfg[322] = { 1'b0, 8'h77, 8'ha8}; // CH=3 OP=1
cfg[323] = { 1'b1, 8'he1, 8'hcd}; // CH=4 OP=0
cfg[324] = { 1'b1, 8'h60, 8'h87}; // CH=3 OP=0
cfg[325] = { 1'b0, 8'h76, 8'h8a}; // CH=2 OP=1
cfg[326] = { 1'b1, 8'ha1, 8'h74}; // CH=4 OP=0
cfg[327] = { 1'b0, 8'h83, 8'h2a}; // CH=3 OP=0
cfg[328] = { 1'b1, 8'he4, 8'h1d}; // CH=3 OP=1
cfg[329] = { 1'b0, 8'hcc, 8'h39}; // CH=0 OP=3
cfg[330] = { 1'b0, 8'h5c, 8'h94}; // CH=0 OP=3
cfg[331] = { 1'b0, 8'h5e, 8'h79}; // CH=2 OP=3
cfg[332] = { 1'b1, 8'hd6, 8'h8a}; // CH=5 OP=1
cfg[333] = { 1'b0, 8'hb7, 8'h57}; // CH=3 OP=1
cfg[334] = { 1'b1, 8'h8d, 8'hdf}; // CH=4 OP=3
cfg[335] = { 1'b1, 8'h69, 8'h8e}; // CH=4 OP=2
cfg[336] = { 1'b1, 8'hd1, 8'h2f}; // CH=4 OP=0
cfg[337] = { 1'b0, 8'h54, 8'h57}; // CH=0 OP=1
cfg[338] = { 1'b1, 8'h39, 8'h75}; // CH=4 OP=2
cfg[339] = { 1'b1, 8'h9b, 8'hae}; // CH=6 OP=2
cfg[340] = { 1'b1, 8'h84, 8'h61}; // CH=3 OP=1
cfg[341] = { 1'b0, 8'h47, 8'hc0}; // CH=3 OP=1
cfg[342] = { 1'b0, 8'h9e, 8'hf3}; // CH=2 OP=3
cfg[343] = { 1'b1, 8'h7d, 8'hc}; // CH=4 OP=3
cfg[344] = { 1'b1, 8'he6, 8'h99}; // CH=5 OP=1
cfg[345] = { 1'b1, 8'hc4, 8'h2}; // CH=3 OP=1
cfg[346] = { 1'b0, 8'hcc, 8'hd3}; // CH=0 OP=3
cfg[347] = { 1'b0, 8'h63, 8'h28}; // CH=3 OP=0
cfg[348] = { 1'b1, 8'h34, 8'h61}; // CH=3 OP=1
cfg[349] = { 1'b1, 8'hcf, 8'h66}; // CH=6 OP=3
cfg[350] = { 1'b0, 8'h53, 8'hc7}; // CH=3 OP=0
cfg[351] = { 1'b1, 8'h68, 8'h87}; // CH=3 OP=2
cfg[352] = { 1'b0, 8'h5b, 8'h1d}; // CH=3 OP=2
cfg[353] = { 1'b0, 8'h67, 8'h6b}; // CH=3 OP=1
cfg[354] = { 1'b0, 8'he6, 8'hd0}; // CH=2 OP=1
cfg[355] = { 1'b0, 8'haa, 8'h3}; // CH=2 OP=2
cfg[356] = { 1'b0, 8'h76, 8'hd7}; // CH=2 OP=1
cfg[357] = { 1'b0, 8'hd9, 8'hff}; // CH=1 OP=2
cfg[358] = { 1'b1, 8'hed, 8'h60}; // CH=4 OP=3
cfg[359] = { 1'b0, 8'hcd, 8'hdd}; // CH=1 OP=3
cfg[360] = { 1'b1, 8'h6a, 8'h30}; // CH=5 OP=2
cfg[361] = { 1'b1, 8'h4e, 8'h99}; // CH=5 OP=3
cfg[362] = { 1'b0, 8'hd1, 8'hf4}; // CH=1 OP=0
cfg[363] = { 1'b1, 8'hd1, 8'h5c}; // CH=4 OP=0
cfg[364] = { 1'b0, 8'hb7, 8'h5d}; // CH=3 OP=1
cfg[365] = { 1'b0, 8'h62, 8'h60}; // CH=2 OP=0
cfg[366] = { 1'b0, 8'hd8, 8'h37}; // CH=0 OP=2
cfg[367] = { 1'b1, 8'hb2, 8'h36}; // CH=5 OP=0
cfg[368] = { 1'b0, 8'hbf, 8'h96}; // CH=3 OP=3
cfg[369] = { 1'b1, 8'h9c, 8'h5c}; // CH=3 OP=3
cfg[370] = { 1'b1, 8'hcd, 8'hea}; // CH=4 OP=3
cfg[371] = { 1'b1, 8'h66, 8'hff}; // CH=5 OP=1
cfg[372] = { 1'b0, 8'h5a, 8'h31}; // CH=2 OP=2
cfg[373] = { 1'b1, 8'hb6, 8'hcf}; // CH=5 OP=1
cfg[374] = { 1'b0, 8'h95, 8'h3d}; // CH=1 OP=1
cfg[375] = { 1'b1, 8'hf7, 8'h74}; // CH=6 OP=1
cfg[376] = { 1'b1, 8'hd0, 8'hab}; // CH=3 OP=0
cfg[377] = { 1'b0, 8'h82, 8'he2}; // CH=2 OP=0
cfg[378] = { 1'b1, 8'h41, 8'h78}; // CH=4 OP=0
cfg[379] = { 1'b0, 8'hde, 8'hd5}; // CH=2 OP=3
cfg[380] = { 1'b1, 8'hab, 8'hbf}; // CH=6 OP=2
cfg[381] = { 1'b1, 8'hef, 8'hbe}; // CH=6 OP=3
cfg[382] = { 1'b1, 8'hbe, 8'h38}; // CH=5 OP=3
cfg[383] = { 1'b0, 8'hfb, 8'h16}; // CH=3 OP=2
cfg[384] = { 1'b1, 8'h6a, 8'hab}; // CH=5 OP=2
cfg[385] = { 1'b1, 8'hf2, 8'ha3}; // CH=5 OP=0
cfg[386] = { 1'b1, 8'hf2, 8'h73}; // CH=5 OP=0
cfg[387] = { 1'b1, 8'hbb, 8'hf5}; // CH=6 OP=2
cfg[388] = { 1'b1, 8'h3a, 8'h36}; // CH=5 OP=2
cfg[389] = { 1'b0, 8'h3b, 8'h14}; // CH=3 OP=2
cfg[390] = { 1'b1, 8'hd0, 8'hbf}; // CH=3 OP=0
cfg[391] = { 1'b1, 8'h3c, 8'hf1}; // CH=3 OP=3
cfg[392] = { 1'b1, 8'h5e, 8'haf}; // CH=5 OP=3
cfg[393] = { 1'b1, 8'h93, 8'hab}; // CH=6 OP=0
cfg[394] = { 1'b1, 8'h3d, 8'h15}; // CH=4 OP=3
cfg[395] = { 1'b0, 8'h92, 8'h7}; // CH=2 OP=0
cfg[396] = { 1'b1, 8'hc9, 8'hfa}; // CH=4 OP=2
cfg[397] = { 1'b0, 8'h78, 8'hb5}; // CH=0 OP=2
cfg[398] = { 1'b0, 8'hfd, 8'hef}; // CH=1 OP=3
cfg[399] = { 1'b1, 8'h40, 8'h2b}; // CH=3 OP=0
cfg[400] = { 1'b0, 8'h42, 8'h55}; // CH=2 OP=0
cfg[401] = { 1'b1, 8'h33, 8'hab}; // CH=6 OP=0
cfg[402] = { 1'b1, 8'he2, 8'h38}; // CH=5 OP=0
cfg[403] = { 1'b1, 8'h8d, 8'hdc}; // CH=4 OP=3
cfg[404] = { 1'b0, 8'ha3, 8'h2b}; // CH=3 OP=0
cfg[405] = { 1'b1, 8'haa, 8'h1d}; // CH=5 OP=2
cfg[406] = { 1'b1, 8'ha4, 8'h82}; // CH=3 OP=1
cfg[407] = { 1'b0, 8'h5a, 8'hdc}; // CH=2 OP=2
cfg[408] = { 1'b1, 8'h49, 8'h6c}; // CH=4 OP=2
cfg[409] = { 1'b0, 8'h74, 8'h11}; // CH=0 OP=1
cfg[410] = { 1'b0, 8'hca, 8'h76}; // CH=2 OP=2
cfg[411] = { 1'b0, 8'h75, 8'hab}; // CH=1 OP=1
cfg[412] = { 1'b1, 8'had, 8'h1c}; // CH=4 OP=3
cfg[413] = { 1'b0, 8'h89, 8'heb}; // CH=1 OP=2
cfg[414] = { 1'b1, 8'hb4, 8'h4d}; // CH=3 OP=1
cfg[415] = { 1'b0, 8'hd1, 8'hed}; // CH=1 OP=0
cfg[416] = { 1'b1, 8'h53, 8'h1e}; // CH=6 OP=0
cfg[417] = { 1'b1, 8'he1, 8'h19}; // CH=4 OP=0
cfg[418] = { 1'b0, 8'hfc, 8'h9c}; // CH=0 OP=3
cfg[419] = { 1'b1, 8'hac, 8'h9f}; // CH=3 OP=3
cfg[420] = { 1'b1, 8'h9f, 8'h69}; // CH=6 OP=3
cfg[421] = { 1'b0, 8'hc4, 8'hde}; // CH=0 OP=1
cfg[422] = { 1'b0, 8'hcc, 8'h8c}; // CH=0 OP=3
cfg[423] = { 1'b1, 8'h62, 8'h15}; // CH=5 OP=0
cfg[424] = { 1'b1, 8'h9a, 8'hca}; // CH=5 OP=2
cfg[425] = { 1'b0, 8'h7d, 8'h9b}; // CH=1 OP=3
cfg[426] = { 1'b0, 8'h47, 8'hef}; // CH=3 OP=1
cfg[427] = { 1'b0, 8'hd3, 8'he6}; // CH=3 OP=0
cfg[428] = { 1'b0, 8'hcf, 8'h11}; // CH=3 OP=3
cfg[429] = { 1'b0, 8'h7c, 8'hb1}; // CH=0 OP=3
cfg[430] = { 1'b1, 8'h5a, 8'h1a}; // CH=5 OP=2
cfg[431] = { 1'b1, 8'h44, 8'hdf}; // CH=3 OP=1
cfg[432] = { 1'b1, 8'h9a, 8'hac}; // CH=5 OP=2
cfg[433] = { 1'b0, 8'h64, 8'h3d}; // CH=0 OP=1
cfg[434] = { 1'b0, 8'h7b, 8'h4d}; // CH=3 OP=2
cfg[435] = { 1'b1, 8'hc3, 8'h2b}; // CH=6 OP=0
cfg[436] = { 1'b1, 8'h96, 8'h11}; // CH=5 OP=1
cfg[437] = { 1'b0, 8'h66, 8'h23}; // CH=2 OP=1
cfg[438] = { 1'b0, 8'he2, 8'hd4}; // CH=2 OP=0
cfg[439] = { 1'b1, 8'hfd, 8'hee}; // CH=4 OP=3
cfg[440] = { 1'b1, 8'hdc, 8'he7}; // CH=3 OP=3
cfg[441] = { 1'b0, 8'h88, 8'h6c}; // CH=0 OP=2
cfg[442] = { 1'b0, 8'h96, 8'h7}; // CH=2 OP=1
cfg[443] = { 1'b1, 8'h3f, 8'h6b}; // CH=6 OP=3
cfg[444] = { 1'b0, 8'h65, 8'h6b}; // CH=1 OP=1
cfg[445] = { 1'b1, 8'h90, 8'h5a}; // CH=3 OP=0
cfg[446] = { 1'b0, 8'ha1, 8'h68}; // CH=1 OP=0
cfg[447] = { 1'b1, 8'hc4, 8'h30}; // CH=3 OP=1
cfg[448] = { 1'b1, 8'h98, 8'h60}; // CH=3 OP=2
cfg[449] = { 1'b1, 8'h87, 8'h1b}; // CH=6 OP=1
cfg[450] = { 1'b0, 8'h6e, 8'h31}; // CH=2 OP=3
cfg[451] = { 1'b0, 8'hdb, 8'h8b}; // CH=3 OP=2
cfg[452] = { 1'b1, 8'he2, 8'hff}; // CH=5 OP=0
cfg[453] = { 1'b1, 8'h4d, 8'hb0}; // CH=4 OP=3
cfg[454] = { 1'b0, 8'hb9, 8'hae}; // CH=1 OP=2
cfg[455] = { 1'b1, 8'h47, 8'h27}; // CH=6 OP=1
cfg[456] = { 1'b0, 8'he9, 8'h7b}; // CH=1 OP=2
cfg[457] = { 1'b1, 8'had, 8'hab}; // CH=4 OP=3
cfg[458] = { 1'b0, 8'h46, 8'hb}; // CH=2 OP=1
cfg[459] = { 1'b1, 8'hcd, 8'h27}; // CH=4 OP=3
cfg[460] = { 1'b1, 8'h3b, 8'h58}; // CH=6 OP=2
cfg[461] = { 1'b1, 8'he2, 8'he3}; // CH=5 OP=0
cfg[462] = { 1'b0, 8'h92, 8'h28}; // CH=2 OP=0
cfg[463] = { 1'b0, 8'h40, 8'h7a}; // CH=0 OP=0
cfg[464] = { 1'b1, 8'h67, 8'h32}; // CH=6 OP=1
cfg[465] = { 1'b0, 8'hcb, 8'h79}; // CH=3 OP=2
cfg[466] = { 1'b0, 8'h39, 8'h62}; // CH=1 OP=2
cfg[467] = { 1'b0, 8'h45, 8'h72}; // CH=1 OP=1
cfg[468] = { 1'b0, 8'h6c, 8'hfd}; // CH=0 OP=3
cfg[469] = { 1'b1, 8'hc4, 8'ha0}; // CH=3 OP=1
cfg[470] = { 1'b0, 8'ha7, 8'h38}; // CH=3 OP=1
cfg[471] = { 1'b1, 8'h89, 8'h4c}; // CH=4 OP=2
cfg[472] = { 1'b1, 8'hb3, 8'h74}; // CH=6 OP=0
cfg[473] = { 1'b1, 8'hb2, 8'h5b}; // CH=5 OP=0
cfg[474] = { 1'b1, 8'hc5, 8'hc2}; // CH=4 OP=1
cfg[475] = { 1'b0, 8'h53, 8'h8e}; // CH=3 OP=0
cfg[476] = { 1'b1, 8'h8c, 8'h90}; // CH=3 OP=3
cfg[477] = { 1'b1, 8'hd1, 8'h3}; // CH=4 OP=0
cfg[478] = { 1'b1, 8'h3d, 8'h0}; // CH=4 OP=3
cfg[479] = { 1'b0, 8'he4, 8'ha1}; // CH=0 OP=1
cfg[480] = { 1'b1, 8'h59, 8'ha8}; // CH=4 OP=2
cfg[481] = { 1'b1, 8'hc7, 8'h31}; // CH=6 OP=1
cfg[482] = { 1'b0, 8'h7a, 8'h4c}; // CH=2 OP=2
cfg[483] = { 1'b1, 8'haa, 8'ha7}; // CH=5 OP=2
cfg[484] = { 1'b0, 8'h44, 8'hf2}; // CH=0 OP=1
cfg[485] = { 1'b0, 8'h41, 8'h45}; // CH=1 OP=0
cfg[486] = { 1'b0, 8'h4e, 8'hd1}; // CH=2 OP=3
cfg[487] = { 1'b1, 8'hb1, 8'ha3}; // CH=4 OP=0
cfg[488] = { 1'b0, 8'h37, 8'he0}; // CH=3 OP=1
cfg[489] = { 1'b1, 8'h8a, 8'he2}; // CH=5 OP=2
cfg[490] = { 1'b1, 8'hbc, 8'h2b}; // CH=3 OP=3
cfg[491] = { 1'b0, 8'hb7, 8'hc5}; // CH=3 OP=1
cfg[492] = { 1'b0, 8'he4, 8'hb0}; // CH=0 OP=1
cfg[493] = { 1'b0, 8'hd6, 8'h1a}; // CH=2 OP=1
cfg[494] = { 1'b1, 8'h7e, 8'h12}; // CH=5 OP=3
cfg[495] = { 1'b0, 8'hcd, 8'hec}; // CH=1 OP=3
cfg[496] = { 1'b0, 8'h7e, 8'h8f}; // CH=2 OP=3
cfg[497] = { 1'b0, 8'hb6, 8'h70}; // CH=2 OP=1
cfg[498] = { 1'b1, 8'hd2, 8'h52}; // CH=5 OP=0
cfg[499] = { 1'b1, 8'h47, 8'hdc}; // CH=6 OP=1
cfg[500] = { 1'b0, 8'h84, 8'h98}; // CH=0 OP=1
cfg[501] = { 1'b0, 8'h3b, 8'ha1}; // CH=3 OP=2
cfg[502] = { 1'b0, 8'h6b, 8'h51}; // CH=3 OP=2
cfg[503] = { 1'b1, 8'h7d, 8'h5a}; // CH=4 OP=3
cfg[504] = { 1'b0, 8'hfc, 8'hd8}; // CH=0 OP=3
cfg[505] = { 1'b1, 8'h8c, 8'h3d}; // CH=3 OP=3
cfg[506] = { 1'b0, 8'hfc, 8'hef}; // CH=0 OP=3
cfg[507] = { 1'b0, 8'h4e, 8'hce}; // CH=2 OP=3
cfg[508] = { 1'b0, 8'hf3, 8'hb3}; // CH=3 OP=0
cfg[509] = { 1'b0, 8'h77, 8'hc3}; // CH=3 OP=1
cfg[510] = { 1'b0, 8'hb2, 8'h64}; // CH=2 OP=0
cfg[511] = { 1'b0, 8'hd1, 8'hb5}; // CH=1 OP=0
cfg[512] = { 1'b1, 8'hc6, 8'h20}; // CH=5 OP=1
cfg[513] = { 1'b1, 8'hd6, 8'h9d}; // CH=5 OP=1
cfg[514] = { 1'b0, 8'hd3, 8'hb4}; // CH=3 OP=0
cfg[515] = { 1'b1, 8'h5f, 8'hf2}; // CH=6 OP=3
cfg[516] = { 1'b1, 8'h5b, 8'he1}; // CH=6 OP=2
cfg[517] = { 1'b1, 8'ha9, 8'hb0}; // CH=4 OP=2
cfg[518] = { 1'b1, 8'hd3, 8'h63}; // CH=6 OP=0
cfg[519] = { 1'b1, 8'h96, 8'h27}; // CH=5 OP=1
cfg[520] = { 1'b0, 8'hfa, 8'hc1}; // CH=2 OP=2
cfg[521] = { 1'b1, 8'haf, 8'h80}; // CH=6 OP=3
cfg[522] = { 1'b0, 8'hcf, 8'h5b}; // CH=3 OP=3
cfg[523] = { 1'b1, 8'h6c, 8'h91}; // CH=3 OP=3
cfg[524] = { 1'b1, 8'hbc, 8'h9f}; // CH=3 OP=3
cfg[525] = { 1'b0, 8'hf4, 8'h13}; // CH=0 OP=1
cfg[526] = { 1'b0, 8'ha4, 8'hdb}; // CH=0 OP=1
cfg[527] = { 1'b1, 8'hf3, 8'h39}; // CH=6 OP=0
cfg[528] = { 1'b0, 8'h89, 8'h2f}; // CH=1 OP=2
cfg[529] = { 1'b0, 8'h84, 8'hf1}; // CH=0 OP=1
cfg[530] = { 1'b1, 8'h33, 8'h71}; // CH=6 OP=0
cfg[531] = { 1'b0, 8'h5d, 8'hcc}; // CH=1 OP=3
cfg[532] = { 1'b1, 8'hfc, 8'h16}; // CH=3 OP=3
cfg[533] = { 1'b0, 8'h4f, 8'hd3}; // CH=3 OP=3
cfg[534] = { 1'b1, 8'h79, 8'hee}; // CH=4 OP=2
cfg[535] = { 1'b0, 8'h54, 8'h65}; // CH=0 OP=1
cfg[536] = { 1'b0, 8'h8d, 8'h84}; // CH=1 OP=3
cfg[537] = { 1'b0, 8'h74, 8'h77}; // CH=0 OP=1
cfg[538] = { 1'b1, 8'h65, 8'h6a}; // CH=4 OP=1
cfg[539] = { 1'b1, 8'hd6, 8'h37}; // CH=5 OP=1
cfg[540] = { 1'b0, 8'ha2, 8'h51}; // CH=2 OP=0
cfg[541] = { 1'b1, 8'h95, 8'h7e}; // CH=4 OP=1
cfg[542] = { 1'b0, 8'h68, 8'hbb}; // CH=0 OP=2
cfg[543] = { 1'b1, 8'h56, 8'h5f}; // CH=5 OP=1
cfg[544] = { 1'b0, 8'hbb, 8'hf7}; // CH=3 OP=2
cfg[545] = { 1'b1, 8'h40, 8'h33}; // CH=3 OP=0
cfg[546] = { 1'b0, 8'hb7, 8'h78}; // CH=3 OP=1
cfg[547] = { 1'b0, 8'hb8, 8'hec}; // CH=0 OP=2
cfg[548] = { 1'b0, 8'h3d, 8'h51}; // CH=1 OP=3
cfg[549] = { 1'b1, 8'hf6, 8'h27}; // CH=5 OP=1
cfg[550] = { 1'b1, 8'hb1, 8'hc9}; // CH=4 OP=0
cfg[551] = { 1'b1, 8'hdc, 8'hc9}; // CH=3 OP=3
cfg[552] = { 1'b0, 8'h98, 8'hc6}; // CH=0 OP=2
cfg[553] = { 1'b0, 8'hf7, 8'h11}; // CH=3 OP=1
cfg[554] = { 1'b1, 8'hee, 8'hd6}; // CH=5 OP=3
cfg[555] = { 1'b0, 8'h7e, 8'hef}; // CH=2 OP=3
cfg[556] = { 1'b1, 8'h36, 8'h99}; // CH=5 OP=1
cfg[557] = { 1'b1, 8'hee, 8'h85}; // CH=5 OP=3
cfg[558] = { 1'b1, 8'hdb, 8'hd6}; // CH=6 OP=2
cfg[559] = { 1'b1, 8'h8c, 8'h22}; // CH=3 OP=3
cfg[560] = { 1'b1, 8'hbb, 8'hd3}; // CH=6 OP=2
cfg[561] = { 1'b0, 8'h80, 8'hb0}; // CH=0 OP=0
cfg[562] = { 1'b0, 8'hac, 8'h48}; // CH=0 OP=3
cfg[563] = { 1'b0, 8'h3e, 8'h3f}; // CH=2 OP=3
cfg[564] = { 1'b1, 8'h4e, 8'h6e}; // CH=5 OP=3
cfg[565] = { 1'b0, 8'he8, 8'hc2}; // CH=0 OP=2
cfg[566] = { 1'b0, 8'h6d, 8'h16}; // CH=1 OP=3
cfg[567] = { 1'b1, 8'h44, 8'h91}; // CH=3 OP=1
cfg[568] = { 1'b1, 8'h41, 8'h6c}; // CH=4 OP=0
cfg[569] = { 1'b1, 8'h32, 8'hf8}; // CH=5 OP=0
cfg[570] = { 1'b0, 8'he2, 8'h99}; // CH=2 OP=0
cfg[571] = { 1'b0, 8'he0, 8'hef}; // CH=0 OP=0
cfg[572] = { 1'b1, 8'h95, 8'h69}; // CH=4 OP=1
cfg[573] = { 1'b0, 8'hc2, 8'h7e}; // CH=2 OP=0
cfg[574] = { 1'b1, 8'h85, 8'h6a}; // CH=4 OP=1
cfg[575] = { 1'b1, 8'h9b, 8'h8d}; // CH=6 OP=2
cfg[576] = { 1'b0, 8'h7e, 8'h9e}; // CH=2 OP=3
cfg[577] = { 1'b1, 8'hc0, 8'h99}; // CH=3 OP=0
cfg[578] = { 1'b0, 8'hc8, 8'h91}; // CH=0 OP=2
cfg[579] = { 1'b0, 8'h61, 8'h45}; // CH=1 OP=0
cfg[580] = { 1'b1, 8'h51, 8'h79}; // CH=4 OP=0
cfg[581] = { 1'b1, 8'ha8, 8'h5a}; // CH=3 OP=2
cfg[582] = { 1'b1, 8'h3e, 8'h6a}; // CH=5 OP=3
cfg[583] = { 1'b1, 8'h5e, 8'he8}; // CH=5 OP=3
cfg[584] = { 1'b0, 8'hdf, 8'h85}; // CH=3 OP=3
cfg[585] = { 1'b0, 8'h7d, 8'h66}; // CH=1 OP=3
cfg[586] = { 1'b1, 8'h58, 8'he4}; // CH=3 OP=2
cfg[587] = { 1'b0, 8'h92, 8'ha4}; // CH=2 OP=0
cfg[588] = { 1'b1, 8'hff, 8'h6d}; // CH=6 OP=3
cfg[589] = { 1'b1, 8'h4e, 8'hce}; // CH=5 OP=3
cfg[590] = { 1'b0, 8'hc7, 8'h1f}; // CH=3 OP=1
cfg[591] = { 1'b0, 8'haa, 8'hc8}; // CH=2 OP=2
cfg[592] = { 1'b0, 8'he2, 8'h6}; // CH=2 OP=0
cfg[593] = { 1'b0, 8'h35, 8'h82}; // CH=1 OP=1
cfg[594] = { 1'b0, 8'hac, 8'hae}; // CH=0 OP=3
cfg[595] = { 1'b0, 8'hf9, 8'h92}; // CH=1 OP=2
cfg[596] = { 1'b0, 8'hdf, 8'hea}; // CH=3 OP=3
cfg[597] = { 1'b1, 8'h57, 8'h7d}; // CH=6 OP=1
cfg[598] = { 1'b0, 8'hd8, 8'h7c}; // CH=0 OP=2
cfg[599] = { 1'b0, 8'hf8, 8'h4a}; // CH=0 OP=2
cfg[600] = { 1'b1, 8'hc0, 8'hdb}; // CH=3 OP=0
cfg[601] = { 1'b0, 8'hc6, 8'hd5}; // CH=2 OP=1
cfg[602] = { 1'b0, 8'hcc, 8'hb8}; // CH=0 OP=3
cfg[603] = { 1'b0, 8'h58, 8'hed}; // CH=0 OP=2
cfg[604] = { 1'b0, 8'ha4, 8'h1}; // CH=0 OP=1
cfg[605] = { 1'b1, 8'h9d, 8'hfe}; // CH=4 OP=3
cfg[606] = { 1'b0, 8'h3a, 8'hde}; // CH=2 OP=2
cfg[607] = { 1'b1, 8'h44, 8'h35}; // CH=3 OP=1
cfg[608] = { 1'b1, 8'h41, 8'h49}; // CH=4 OP=0
cfg[609] = { 1'b1, 8'hd2, 8'h14}; // CH=5 OP=0
cfg[610] = { 1'b0, 8'h44, 8'hd4}; // CH=0 OP=1
cfg[611] = { 1'b0, 8'hfc, 8'h6e}; // CH=0 OP=3
cfg[612] = { 1'b1, 8'he9, 8'h51}; // CH=4 OP=2
cfg[613] = { 1'b1, 8'hea, 8'he1}; // CH=5 OP=2
cfg[614] = { 1'b0, 8'h7e, 8'h86}; // CH=2 OP=3
cfg[615] = { 1'b1, 8'hfc, 8'h23}; // CH=3 OP=3
cfg[616] = { 1'b1, 8'hf7, 8'h5d}; // CH=6 OP=1
cfg[617] = { 1'b0, 8'h6e, 8'ha1}; // CH=2 OP=3
cfg[618] = { 1'b1, 8'haf, 8'hbd}; // CH=6 OP=3
cfg[619] = { 1'b0, 8'h81, 8'hd2}; // CH=1 OP=0
cfg[620] = { 1'b1, 8'h90, 8'ha6}; // CH=3 OP=0
cfg[621] = { 1'b1, 8'hfe, 8'h41}; // CH=5 OP=3
cfg[622] = { 1'b1, 8'h4f, 8'ha8}; // CH=6 OP=3
cfg[623] = { 1'b0, 8'h31, 8'h67}; // CH=1 OP=0
cfg[624] = { 1'b0, 8'hb7, 8'h2c}; // CH=3 OP=1
cfg[625] = { 1'b0, 8'hda, 8'hef}; // CH=2 OP=2
cfg[626] = { 1'b0, 8'h37, 8'h90}; // CH=3 OP=1
cfg[627] = { 1'b1, 8'hd8, 8'h66}; // CH=3 OP=2
cfg[628] = { 1'b1, 8'h95, 8'h85}; // CH=4 OP=1
cfg[629] = { 1'b0, 8'h67, 8'h37}; // CH=3 OP=1
cfg[630] = { 1'b0, 8'hd4, 8'h58}; // CH=0 OP=1
cfg[631] = { 1'b1, 8'hd2, 8'h4f}; // CH=5 OP=0
cfg[632] = { 1'b0, 8'h68, 8'hf7}; // CH=0 OP=2
cfg[633] = { 1'b0, 8'h9d, 8'h53}; // CH=1 OP=3
cfg[634] = { 1'b0, 8'h4f, 8'ha}; // CH=3 OP=3
cfg[635] = { 1'b1, 8'hfe, 8'he4}; // CH=5 OP=3
cfg[636] = { 1'b1, 8'ha3, 8'h1b}; // CH=6 OP=0
cfg[637] = { 1'b1, 8'hb7, 8'hf3}; // CH=6 OP=1
cfg[638] = { 1'b0, 8'h79, 8'h88}; // CH=1 OP=2
cfg[639] = { 1'b0, 8'hbd, 8'hf0}; // CH=1 OP=3
cfg[640] = { 1'b0, 8'h91, 8'hfe}; // CH=1 OP=0
cfg[641] = { 1'b0, 8'h64, 8'h4d}; // CH=0 OP=1
cfg[642] = { 1'b0, 8'h86, 8'h44}; // CH=2 OP=1
cfg[643] = { 1'b1, 8'hd9, 8'ha2}; // CH=4 OP=2
cfg[644] = { 1'b0, 8'he3, 8'h2d}; // CH=3 OP=0
cfg[645] = { 1'b1, 8'hc7, 8'ha6}; // CH=6 OP=1
cfg[646] = { 1'b1, 8'he2, 8'hb0}; // CH=5 OP=0
cfg[647] = { 1'b1, 8'hd5, 8'h1f}; // CH=4 OP=1
cfg[648] = { 1'b0, 8'h5d, 8'h14}; // CH=1 OP=3
cfg[649] = { 1'b1, 8'h4d, 8'h40}; // CH=4 OP=3
cfg[650] = { 1'b1, 8'h4b, 8'hc4}; // CH=6 OP=2
cfg[651] = { 1'b0, 8'h98, 8'h6}; // CH=0 OP=2
cfg[652] = { 1'b0, 8'hdc, 8'h67}; // CH=0 OP=3
cfg[653] = { 1'b0, 8'h7f, 8'h30}; // CH=3 OP=3
cfg[654] = { 1'b1, 8'hac, 8'h96}; // CH=3 OP=3
cfg[655] = { 1'b0, 8'h52, 8'h4b}; // CH=2 OP=0
cfg[656] = { 1'b1, 8'h56, 8'hff}; // CH=5 OP=1
cfg[657] = { 1'b0, 8'h64, 8'hfa}; // CH=0 OP=1
cfg[658] = { 1'b0, 8'heb, 8'h58}; // CH=3 OP=2
cfg[659] = { 1'b0, 8'h30, 8'ha5}; // CH=0 OP=0
cfg[660] = { 1'b0, 8'h41, 8'hf1}; // CH=1 OP=0
cfg[661] = { 1'b1, 8'ha8, 8'h41}; // CH=3 OP=2
cfg[662] = { 1'b0, 8'hd8, 8'h2}; // CH=0 OP=2
cfg[663] = { 1'b1, 8'h6e, 8'h9b}; // CH=5 OP=3
cfg[664] = { 1'b1, 8'hb9, 8'h18}; // CH=4 OP=2
cfg[665] = { 1'b1, 8'hb8, 8'h5b}; // CH=3 OP=2
cfg[666] = { 1'b0, 8'h7b, 8'h81}; // CH=3 OP=2
cfg[667] = { 1'b0, 8'hd3, 8'h3e}; // CH=3 OP=0
cfg[668] = { 1'b0, 8'h79, 8'hb4}; // CH=1 OP=2
cfg[669] = { 1'b0, 8'h6a, 8'hee}; // CH=2 OP=2
cfg[670] = { 1'b1, 8'hf3, 8'h2f}; // CH=6 OP=0
cfg[671] = { 1'b1, 8'h59, 8'hd7}; // CH=4 OP=2
cfg[672] = { 1'b1, 8'h3e, 8'haf}; // CH=5 OP=3
cfg[673] = { 1'b0, 8'hcf, 8'h1d}; // CH=3 OP=3
cfg[674] = { 1'b0, 8'hb3, 8'hd7}; // CH=3 OP=0
cfg[675] = { 1'b0, 8'h99, 8'h8f}; // CH=1 OP=2
cfg[676] = { 1'b1, 8'ha1, 8'h9e}; // CH=4 OP=0
cfg[677] = { 1'b0, 8'hdf, 8'h10}; // CH=3 OP=3
cfg[678] = { 1'b0, 8'h93, 8'h6e}; // CH=3 OP=0
cfg[679] = { 1'b1, 8'h81, 8'hfd}; // CH=4 OP=0
cfg[680] = { 1'b1, 8'hb1, 8'h92}; // CH=4 OP=0
cfg[681] = { 1'b0, 8'h88, 8'h69}; // CH=0 OP=2
cfg[682] = { 1'b0, 8'h38, 8'h42}; // CH=0 OP=2
cfg[683] = { 1'b0, 8'h55, 8'hb7}; // CH=1 OP=1
cfg[684] = { 1'b0, 8'ha9, 8'h43}; // CH=1 OP=2
cfg[685] = { 1'b1, 8'h42, 8'hbc}; // CH=5 OP=0
cfg[686] = { 1'b0, 8'he3, 8'h5a}; // CH=3 OP=0
cfg[687] = { 1'b1, 8'hc2, 8'h6a}; // CH=5 OP=0
cfg[688] = { 1'b1, 8'h55, 8'hd9}; // CH=4 OP=1
cfg[689] = { 1'b0, 8'hd6, 8'hd6}; // CH=2 OP=1
cfg[690] = { 1'b1, 8'h87, 8'h68}; // CH=6 OP=1
cfg[691] = { 1'b1, 8'h73, 8'hd2}; // CH=6 OP=0
cfg[692] = { 1'b0, 8'h9a, 8'h48}; // CH=2 OP=2
cfg[693] = { 1'b1, 8'h90, 8'h9d}; // CH=3 OP=0
cfg[694] = { 1'b1, 8'h39, 8'hca}; // CH=4 OP=2
cfg[695] = { 1'b0, 8'h7b, 8'h86}; // CH=3 OP=2
cfg[696] = { 1'b1, 8'h5e, 8'he0}; // CH=5 OP=3
cfg[697] = { 1'b0, 8'h79, 8'h4a}; // CH=1 OP=2
cfg[698] = { 1'b1, 8'hdb, 8'h75}; // CH=6 OP=2
cfg[699] = { 1'b1, 8'hd8, 8'h4b}; // CH=3 OP=2
cfg[700] = { 1'b0, 8'h63, 8'hd3}; // CH=3 OP=0
cfg[701] = { 1'b0, 8'hd7, 8'he3}; // CH=3 OP=1
cfg[702] = { 1'b0, 8'h71, 8'h2b}; // CH=1 OP=0
cfg[703] = { 1'b0, 8'h92, 8'hc8}; // CH=2 OP=0
cfg[704] = { 1'b0, 8'hb5, 8'h5d}; // CH=1 OP=1
cfg[705] = { 1'b0, 8'h74, 8'hf8}; // CH=0 OP=1
cfg[706] = { 1'b1, 8'hed, 8'h33}; // CH=4 OP=3
cfg[707] = { 1'b0, 8'hc8, 8'ha8}; // CH=0 OP=2
cfg[708] = { 1'b0, 8'ha0, 8'hf3}; // CH=0 OP=0
cfg[709] = { 1'b0, 8'hf6, 8'hc6}; // CH=2 OP=1
cfg[710] = { 1'b1, 8'h3e, 8'hdb}; // CH=5 OP=3
cfg[711] = { 1'b0, 8'h52, 8'h4c}; // CH=2 OP=0
cfg[712] = { 1'b1, 8'h75, 8'h4d}; // CH=4 OP=1
cfg[713] = { 1'b1, 8'hd3, 8'h87}; // CH=6 OP=0
cfg[714] = { 1'b0, 8'hff, 8'h3c}; // CH=3 OP=3
cfg[715] = { 1'b0, 8'h74, 8'h4f}; // CH=0 OP=1
cfg[716] = { 1'b1, 8'h61, 8'h82}; // CH=4 OP=0
cfg[717] = { 1'b0, 8'h4a, 8'h2a}; // CH=2 OP=2
cfg[718] = { 1'b1, 8'he4, 8'hca}; // CH=3 OP=1
cfg[719] = { 1'b0, 8'h8d, 8'h2}; // CH=1 OP=3
cfg[720] = { 1'b1, 8'h62, 8'h40}; // CH=5 OP=0
cfg[721] = { 1'b1, 8'hff, 8'h93}; // CH=6 OP=3
cfg[722] = { 1'b0, 8'hc9, 8'h8}; // CH=1 OP=2
cfg[723] = { 1'b1, 8'hdb, 8'h76}; // CH=6 OP=2
cfg[724] = { 1'b1, 8'h4f, 8'h54}; // CH=6 OP=3
cfg[725] = { 1'b0, 8'hb0, 8'hd6}; // CH=0 OP=0
cfg[726] = { 1'b0, 8'hda, 8'h0}; // CH=2 OP=2
cfg[727] = { 1'b0, 8'ha5, 8'h1e}; // CH=1 OP=1
cfg[728] = { 1'b0, 8'h73, 8'h2}; // CH=3 OP=0
cfg[729] = { 1'b0, 8'hbd, 8'h8f}; // CH=1 OP=3
cfg[730] = { 1'b1, 8'h50, 8'h12}; // CH=3 OP=0
cfg[731] = { 1'b0, 8'h58, 8'h55}; // CH=0 OP=2
cfg[732] = { 1'b1, 8'h34, 8'h1e}; // CH=3 OP=1
cfg[733] = { 1'b1, 8'h4c, 8'h24}; // CH=3 OP=3
cfg[734] = { 1'b0, 8'h87, 8'h5e}; // CH=3 OP=1
cfg[735] = { 1'b1, 8'hab, 8'he}; // CH=6 OP=2
cfg[736] = { 1'b1, 8'h6d, 8'he9}; // CH=4 OP=3
cfg[737] = { 1'b0, 8'h6f, 8'h94}; // CH=3 OP=3
cfg[738] = { 1'b1, 8'hff, 8'h11}; // CH=6 OP=3
cfg[739] = { 1'b0, 8'hf0, 8'hce}; // CH=0 OP=0
cfg[740] = { 1'b1, 8'he1, 8'h1e}; // CH=4 OP=0
cfg[741] = { 1'b0, 8'ha4, 8'h76}; // CH=0 OP=1
cfg[742] = { 1'b0, 8'hc8, 8'h95}; // CH=0 OP=2
cfg[743] = { 1'b1, 8'h41, 8'he2}; // CH=4 OP=0
cfg[744] = { 1'b1, 8'h90, 8'h69}; // CH=3 OP=0
cfg[745] = { 1'b0, 8'hdf, 8'h14}; // CH=3 OP=3
cfg[746] = { 1'b1, 8'h4d, 8'h2e}; // CH=4 OP=3
cfg[747] = { 1'b1, 8'hbc, 8'hc3}; // CH=3 OP=3
cfg[748] = { 1'b0, 8'hbb, 8'hd4}; // CH=3 OP=2
cfg[749] = { 1'b1, 8'hac, 8'ha2}; // CH=3 OP=3
cfg[750] = { 1'b0, 8'h8d, 8'hc0}; // CH=1 OP=3
cfg[751] = { 1'b0, 8'h8d, 8'h36}; // CH=1 OP=3
cfg[752] = { 1'b0, 8'he1, 8'he1}; // CH=1 OP=0
cfg[753] = { 1'b0, 8'hb2, 8'h4}; // CH=2 OP=0
cfg[754] = { 1'b1, 8'hd8, 8'hb2}; // CH=3 OP=2
cfg[755] = { 1'b0, 8'he7, 8'h91}; // CH=3 OP=1
cfg[756] = { 1'b0, 8'h84, 8'hde}; // CH=0 OP=1
cfg[757] = { 1'b1, 8'h47, 8'h9b}; // CH=6 OP=1
cfg[758] = { 1'b0, 8'he9, 8'hdf}; // CH=1 OP=2
cfg[759] = { 1'b0, 8'ha9, 8'hcd}; // CH=1 OP=2
cfg[760] = { 1'b1, 8'he0, 8'h41}; // CH=3 OP=0
cfg[761] = { 1'b0, 8'hc1, 8'h5a}; // CH=1 OP=0
cfg[762] = { 1'b1, 8'h5b, 8'h3b}; // CH=6 OP=2
cfg[763] = { 1'b1, 8'hb1, 8'h5d}; // CH=4 OP=0
cfg[764] = { 1'b1, 8'h33, 8'he5}; // CH=6 OP=0
cfg[765] = { 1'b0, 8'he3, 8'hcc}; // CH=3 OP=0
cfg[766] = { 1'b1, 8'h57, 8'h50}; // CH=6 OP=1
cfg[767] = { 1'b0, 8'h9e, 8'h73}; // CH=2 OP=3
cfg[768] = { 1'b0, 8'h88, 8'h52}; // CH=0 OP=2
cfg[769] = { 1'b1, 8'h31, 8'h20}; // CH=4 OP=0
cfg[770] = { 1'b0, 8'hbb, 8'h61}; // CH=3 OP=2
cfg[771] = { 1'b0, 8'hf6, 8'h5e}; // CH=2 OP=1
cfg[772] = { 1'b0, 8'h53, 8'ha1}; // CH=3 OP=0
cfg[773] = { 1'b1, 8'h62, 8'h52}; // CH=5 OP=0
cfg[774] = { 1'b1, 8'hed, 8'h85}; // CH=4 OP=3
cfg[775] = { 1'b1, 8'h3e, 8'h82}; // CH=5 OP=3
cfg[776] = { 1'b0, 8'hb1, 8'h9c}; // CH=1 OP=0
cfg[777] = { 1'b0, 8'he6, 8'hc}; // CH=2 OP=1
cfg[778] = { 1'b1, 8'h82, 8'h23}; // CH=5 OP=0
cfg[779] = { 1'b1, 8'ha1, 8'h29}; // CH=4 OP=0
cfg[780] = { 1'b0, 8'hff, 8'hfc}; // CH=3 OP=3
cfg[781] = { 1'b1, 8'ha0, 8'h2a}; // CH=3 OP=0
cfg[782] = { 1'b0, 8'hf3, 8'h65}; // CH=3 OP=0
cfg[783] = { 1'b1, 8'h78, 8'h86}; // CH=3 OP=2
cfg[784] = { 1'b0, 8'he1, 8'h74}; // CH=1 OP=0
cfg[785] = { 1'b0, 8'ha1, 8'hb2}; // CH=1 OP=0
cfg[786] = { 1'b0, 8'h66, 8'h63}; // CH=2 OP=1
cfg[787] = { 1'b0, 8'h8a, 8'h9a}; // CH=2 OP=2
cfg[788] = { 1'b0, 8'hbd, 8'h1c}; // CH=1 OP=3
cfg[789] = { 1'b1, 8'hbc, 8'h24}; // CH=3 OP=3
cfg[790] = { 1'b0, 8'h5c, 8'h4e}; // CH=0 OP=3
cfg[791] = { 1'b1, 8'h4f, 8'hb3}; // CH=6 OP=3
cfg[792] = { 1'b0, 8'hc8, 8'h3a}; // CH=0 OP=2
cfg[793] = { 1'b0, 8'ha9, 8'hae}; // CH=1 OP=2
cfg[794] = { 1'b0, 8'h4b, 8'h60}; // CH=3 OP=2
cfg[795] = { 1'b0, 8'h4b, 8'hc3}; // CH=3 OP=2
cfg[796] = { 1'b0, 8'h31, 8'h29}; // CH=1 OP=0
cfg[797] = { 1'b0, 8'h30, 8'hb3}; // CH=0 OP=0
cfg[798] = { 1'b0, 8'h58, 8'hc2}; // CH=0 OP=2
cfg[799] = { 1'b1, 8'h7c, 8'h12}; // CH=3 OP=3
cfg[800] = { 1'b1, 8'hca, 8'h98}; // CH=5 OP=2
cfg[801] = { 1'b0, 8'h7d, 8'ha9}; // CH=1 OP=3
cfg[802] = { 1'b1, 8'hb7, 8'ha7}; // CH=6 OP=1
cfg[803] = { 1'b1, 8'h65, 8'h95}; // CH=4 OP=1
cfg[804] = { 1'b1, 8'hc5, 8'hf5}; // CH=4 OP=1
cfg[805] = { 1'b0, 8'h88, 8'h63}; // CH=0 OP=2
cfg[806] = { 1'b1, 8'hb2, 8'hec}; // CH=5 OP=0
cfg[807] = { 1'b0, 8'h65, 8'he}; // CH=1 OP=1
cfg[808] = { 1'b0, 8'h48, 8'h4d}; // CH=0 OP=2
cfg[809] = { 1'b0, 8'hd2, 8'ha0}; // CH=2 OP=0
cfg[810] = { 1'b0, 8'h7c, 8'h14}; // CH=0 OP=3
cfg[811] = { 1'b0, 8'h9f, 8'h77}; // CH=3 OP=3
cfg[812] = { 1'b1, 8'h78, 8'hb9}; // CH=3 OP=2
cfg[813] = { 1'b0, 8'h98, 8'hca}; // CH=0 OP=2
cfg[814] = { 1'b0, 8'hfe, 8'h53}; // CH=2 OP=3
cfg[815] = { 1'b1, 8'h6a, 8'h9f}; // CH=5 OP=2
cfg[816] = { 1'b0, 8'h92, 8'h59}; // CH=2 OP=0
cfg[817] = { 1'b0, 8'hcc, 8'ha2}; // CH=0 OP=3
cfg[818] = { 1'b1, 8'h9f, 8'ha2}; // CH=6 OP=3
cfg[819] = { 1'b1, 8'h83, 8'hb6}; // CH=6 OP=0
cfg[820] = { 1'b1, 8'hd0, 8'h3e}; // CH=3 OP=0
cfg[821] = { 1'b1, 8'h48, 8'h28}; // CH=3 OP=2
cfg[822] = { 1'b0, 8'he0, 8'hf2}; // CH=0 OP=0
cfg[823] = { 1'b0, 8'he3, 8'h45}; // CH=3 OP=0
cfg[824] = { 1'b0, 8'h83, 8'h4a}; // CH=3 OP=0
cfg[825] = { 1'b0, 8'hef, 8'hb5}; // CH=3 OP=3
cfg[826] = { 1'b0, 8'h7f, 8'h47}; // CH=3 OP=3
cfg[827] = { 1'b0, 8'hb0, 8'h14}; // CH=0 OP=0
cfg[828] = { 1'b0, 8'h4c, 8'hb3}; // CH=0 OP=3
cfg[829] = { 1'b0, 8'hcf, 8'hce}; // CH=3 OP=3
cfg[830] = { 1'b1, 8'hf2, 8'hc}; // CH=5 OP=0
cfg[831] = { 1'b0, 8'h5c, 8'h4}; // CH=0 OP=3
cfg[832] = { 1'b0, 8'h3d, 8'hd}; // CH=1 OP=3
cfg[833] = { 1'b0, 8'h9d, 8'h52}; // CH=1 OP=3
cfg[834] = { 1'b1, 8'h52, 8'hda}; // CH=5 OP=0
cfg[835] = { 1'b0, 8'h99, 8'hf6}; // CH=1 OP=2
cfg[836] = { 1'b0, 8'had, 8'hb4}; // CH=1 OP=3
cfg[837] = { 1'b0, 8'h60, 8'h14}; // CH=0 OP=0
cfg[838] = { 1'b0, 8'hde, 8'h2a}; // CH=2 OP=3
cfg[839] = { 1'b0, 8'hd0, 8'h3b}; // CH=0 OP=0
cfg[840] = { 1'b0, 8'heb, 8'h3f}; // CH=3 OP=2
cfg[841] = { 1'b0, 8'hf8, 8'he9}; // CH=0 OP=2
cfg[842] = { 1'b1, 8'h4a, 8'h4b}; // CH=5 OP=2
cfg[843] = { 1'b0, 8'he7, 8'h63}; // CH=3 OP=1
cfg[844] = { 1'b1, 8'h39, 8'h3d}; // CH=4 OP=2
cfg[845] = { 1'b0, 8'hd3, 8'h34}; // CH=3 OP=0
cfg[846] = { 1'b0, 8'h80, 8'he8}; // CH=0 OP=0
cfg[847] = { 1'b0, 8'he1, 8'hfd}; // CH=1 OP=0
cfg[848] = { 1'b1, 8'h33, 8'h27}; // CH=6 OP=0
cfg[849] = { 1'b1, 8'h89, 8'h4a}; // CH=4 OP=2
cfg[850] = { 1'b0, 8'h72, 8'hf6}; // CH=2 OP=0
cfg[851] = { 1'b0, 8'hbd, 8'h11}; // CH=1 OP=3
cfg[852] = { 1'b1, 8'h5e, 8'h4d}; // CH=5 OP=3
cfg[853] = { 1'b0, 8'h92, 8'h9f}; // CH=2 OP=0
cfg[854] = { 1'b1, 8'h7a, 8'h23}; // CH=5 OP=2
cfg[855] = { 1'b1, 8'h77, 8'h69}; // CH=6 OP=1
cfg[856] = { 1'b0, 8'h9f, 8'hbe}; // CH=3 OP=3
cfg[857] = { 1'b0, 8'h34, 8'hf1}; // CH=0 OP=1
cfg[858] = { 1'b0, 8'h4c, 8'hf5}; // CH=0 OP=3
cfg[859] = { 1'b0, 8'h42, 8'he3}; // CH=2 OP=0
cfg[860] = { 1'b0, 8'h53, 8'hca}; // CH=3 OP=0
cfg[861] = { 1'b0, 8'ha1, 8'hfb}; // CH=1 OP=0
cfg[862] = { 1'b0, 8'hce, 8'h13}; // CH=2 OP=3
cfg[863] = { 1'b0, 8'h6d, 8'h65}; // CH=1 OP=3
cfg[864] = { 1'b0, 8'h90, 8'h8a}; // CH=0 OP=0
cfg[865] = { 1'b1, 8'hf9, 8'h30}; // CH=4 OP=2
cfg[866] = { 1'b0, 8'hb8, 8'hb6}; // CH=0 OP=2
cfg[867] = { 1'b1, 8'ha9, 8'h4c}; // CH=4 OP=2
cfg[868] = { 1'b0, 8'h9e, 8'h2d}; // CH=2 OP=3
cfg[869] = { 1'b0, 8'h82, 8'h97}; // CH=2 OP=0
cfg[870] = { 1'b0, 8'h4c, 8'h73}; // CH=0 OP=3
cfg[871] = { 1'b1, 8'h47, 8'hd}; // CH=6 OP=1
cfg[872] = { 1'b0, 8'h5a, 8'hc8}; // CH=2 OP=2
cfg[873] = { 1'b0, 8'hc0, 8'he0}; // CH=0 OP=0
cfg[874] = { 1'b1, 8'h4a, 8'h8b}; // CH=5 OP=2
cfg[875] = { 1'b1, 8'h7a, 8'hb0}; // CH=5 OP=2
cfg[876] = { 1'b1, 8'h31, 8'h4c}; // CH=4 OP=0
cfg[877] = { 1'b1, 8'h7d, 8'h88}; // CH=4 OP=3
cfg[878] = { 1'b0, 8'haa, 8'hf8}; // CH=2 OP=2
cfg[879] = { 1'b1, 8'h41, 8'hb4}; // CH=4 OP=0
cfg[880] = { 1'b1, 8'hb5, 8'hb2}; // CH=4 OP=1
cfg[881] = { 1'b1, 8'hc2, 8'h3}; // CH=5 OP=0
cfg[882] = { 1'b0, 8'h8a, 8'hf6}; // CH=2 OP=2
cfg[883] = { 1'b0, 8'h6b, 8'hb6}; // CH=3 OP=2
cfg[884] = { 1'b0, 8'hf6, 8'he4}; // CH=2 OP=1
cfg[885] = { 1'b1, 8'ha6, 8'ha1}; // CH=5 OP=1
cfg[886] = { 1'b1, 8'hf2, 8'h58}; // CH=5 OP=0
cfg[887] = { 1'b0, 8'h7a, 8'hc7}; // CH=2 OP=2
cfg[888] = { 1'b0, 8'h72, 8'he0}; // CH=2 OP=0
cfg[889] = { 1'b0, 8'h46, 8'h97}; // CH=2 OP=1
cfg[890] = { 1'b0, 8'hfb, 8'hd8}; // CH=3 OP=2
cfg[891] = { 1'b1, 8'hbd, 8'hdc}; // CH=4 OP=3
cfg[892] = { 1'b1, 8'h48, 8'hd2}; // CH=3 OP=2
cfg[893] = { 1'b1, 8'hb3, 8'h88}; // CH=6 OP=0
cfg[894] = { 1'b0, 8'ha9, 8'h6c}; // CH=1 OP=2
cfg[895] = { 1'b1, 8'h4f, 8'he}; // CH=6 OP=3
cfg[896] = { 1'b0, 8'h41, 8'h66}; // CH=1 OP=0
cfg[897] = { 1'b1, 8'hbc, 8'h2e}; // CH=3 OP=3
cfg[898] = { 1'b1, 8'h45, 8'he}; // CH=4 OP=1
cfg[899] = { 1'b1, 8'h8b, 8'h55}; // CH=6 OP=2
cfg[900] = { 1'b1, 8'h86, 8'h2d}; // CH=5 OP=1
cfg[901] = { 1'b0, 8'h44, 8'h9}; // CH=0 OP=1
cfg[902] = { 1'b1, 8'h8c, 8'hdb}; // CH=3 OP=3
cfg[903] = { 1'b0, 8'h3f, 8'h64}; // CH=3 OP=3
cfg[904] = { 1'b0, 8'he8, 8'hd0}; // CH=0 OP=2
cfg[905] = { 1'b1, 8'h37, 8'hde}; // CH=6 OP=1
cfg[906] = { 1'b0, 8'h78, 8'h45}; // CH=0 OP=2
cfg[907] = { 1'b1, 8'h34, 8'h73}; // CH=3 OP=1
cfg[908] = { 1'b0, 8'h63, 8'h81}; // CH=3 OP=0
cfg[909] = { 1'b1, 8'hb8, 8'h26}; // CH=3 OP=2
cfg[910] = { 1'b1, 8'he5, 8'h9b}; // CH=4 OP=1
cfg[911] = { 1'b1, 8'hef, 8'h65}; // CH=6 OP=3
cfg[912] = { 1'b1, 8'hca, 8'h50}; // CH=5 OP=2
cfg[913] = { 1'b1, 8'h58, 8'h82}; // CH=3 OP=2
cfg[914] = { 1'b1, 8'h40, 8'hff}; // CH=3 OP=0
cfg[915] = { 1'b0, 8'h77, 8'hdd}; // CH=3 OP=1
cfg[916] = { 1'b0, 8'hf0, 8'h22}; // CH=0 OP=0
cfg[917] = { 1'b1, 8'h87, 8'h95}; // CH=6 OP=1
cfg[918] = { 1'b1, 8'h3f, 8'h3c}; // CH=6 OP=3
cfg[919] = { 1'b0, 8'h53, 8'hd7}; // CH=3 OP=0
cfg[920] = { 1'b0, 8'he1, 8'h14}; // CH=1 OP=0
cfg[921] = { 1'b0, 8'hfa, 8'hde}; // CH=2 OP=2
cfg[922] = { 1'b1, 8'h53, 8'hd}; // CH=6 OP=0
cfg[923] = { 1'b0, 8'h93, 8'hc}; // CH=3 OP=0
cfg[924] = { 1'b0, 8'hfb, 8'he9}; // CH=3 OP=2
cfg[925] = { 1'b0, 8'hb8, 8'ha1}; // CH=0 OP=2
cfg[926] = { 1'b1, 8'hf4, 8'h75}; // CH=3 OP=1
cfg[927] = { 1'b0, 8'hcc, 8'h7f}; // CH=0 OP=3
cfg[928] = { 1'b1, 8'hb3, 8'hd2}; // CH=6 OP=0
cfg[929] = { 1'b1, 8'hae, 8'hfe}; // CH=5 OP=3
cfg[930] = { 1'b0, 8'h96, 8'hb}; // CH=2 OP=1
cfg[931] = { 1'b1, 8'h9f, 8'h94}; // CH=6 OP=3
cfg[932] = { 1'b1, 8'h9a, 8'hc}; // CH=5 OP=2
cfg[933] = { 1'b0, 8'hba, 8'hae}; // CH=2 OP=2
cfg[934] = { 1'b0, 8'h61, 8'h66}; // CH=1 OP=0
cfg[935] = { 1'b1, 8'h47, 8'h5a}; // CH=6 OP=1
cfg[936] = { 1'b0, 8'h53, 8'h26}; // CH=3 OP=0
cfg[937] = { 1'b0, 8'h72, 8'h2f}; // CH=2 OP=0
cfg[938] = { 1'b0, 8'h70, 8'hc4}; // CH=0 OP=0
cfg[939] = { 1'b0, 8'h7b, 8'h68}; // CH=3 OP=2
cfg[940] = { 1'b1, 8'h92, 8'hfe}; // CH=5 OP=0
cfg[941] = { 1'b1, 8'h93, 8'h28}; // CH=6 OP=0
cfg[942] = { 1'b1, 8'h9f, 8'h54}; // CH=6 OP=3
cfg[943] = { 1'b1, 8'h4d, 8'h9e}; // CH=4 OP=3
cfg[944] = { 1'b1, 8'hb3, 8'h16}; // CH=6 OP=0
cfg[945] = { 1'b0, 8'hd2, 8'h3}; // CH=2 OP=0
cfg[946] = { 1'b1, 8'had, 8'h34}; // CH=4 OP=3
cfg[947] = { 1'b1, 8'h9f, 8'h97}; // CH=6 OP=3
cfg[948] = { 1'b1, 8'h3f, 8'h8}; // CH=6 OP=3
cfg[949] = { 1'b1, 8'he0, 8'h83}; // CH=3 OP=0
cfg[950] = { 1'b1, 8'hb6, 8'h16}; // CH=5 OP=1
cfg[951] = { 1'b1, 8'h48, 8'heb}; // CH=3 OP=2
cfg[952] = { 1'b0, 8'h96, 8'ha8}; // CH=2 OP=1
cfg[953] = { 1'b0, 8'h49, 8'hbe}; // CH=1 OP=2
cfg[954] = { 1'b0, 8'h57, 8'hc1}; // CH=3 OP=1
cfg[955] = { 1'b0, 8'h8c, 8'h30}; // CH=0 OP=3
cfg[956] = { 1'b1, 8'hef, 8'hdd}; // CH=6 OP=3
cfg[957] = { 1'b1, 8'ha5, 8'h7d}; // CH=4 OP=1
cfg[958] = { 1'b0, 8'h9d, 8'ha6}; // CH=1 OP=3
cfg[959] = { 1'b0, 8'hb3, 8'h3e}; // CH=3 OP=0
cfg[960] = { 1'b0, 8'h9e, 8'he7}; // CH=2 OP=3
cfg[961] = { 1'b0, 8'hf8, 8'h30}; // CH=0 OP=2
cfg[962] = { 1'b0, 8'h7c, 8'hc6}; // CH=0 OP=3
cfg[963] = { 1'b0, 8'h8b, 8'hf}; // CH=3 OP=2
cfg[964] = { 1'b1, 8'h6b, 8'h67}; // CH=6 OP=2
cfg[965] = { 1'b1, 8'h71, 8'hf3}; // CH=4 OP=0
cfg[966] = { 1'b0, 8'ha5, 8'he2}; // CH=1 OP=1
cfg[967] = { 1'b1, 8'h62, 8'hb3}; // CH=5 OP=0
cfg[968] = { 1'b0, 8'hff, 8'hdb}; // CH=3 OP=3
cfg[969] = { 1'b0, 8'hb2, 8'h1a}; // CH=2 OP=0
cfg[970] = { 1'b0, 8'h50, 8'h1}; // CH=0 OP=0
cfg[971] = { 1'b0, 8'h48, 8'h31}; // CH=0 OP=2
cfg[972] = { 1'b0, 8'hc5, 8'hf7}; // CH=1 OP=1
cfg[973] = { 1'b0, 8'h50, 8'h7}; // CH=0 OP=0
cfg[974] = { 1'b1, 8'hbb, 8'h6e}; // CH=6 OP=2
cfg[975] = { 1'b0, 8'h36, 8'h61}; // CH=2 OP=1
cfg[976] = { 1'b1, 8'hdc, 8'h3a}; // CH=3 OP=3
cfg[977] = { 1'b1, 8'h3e, 8'hed}; // CH=5 OP=3
cfg[978] = { 1'b1, 8'h3d, 8'hc9}; // CH=4 OP=3
cfg[979] = { 1'b1, 8'hef, 8'he3}; // CH=6 OP=3
cfg[980] = { 1'b1, 8'h3f, 8'he4}; // CH=6 OP=3
cfg[981] = { 1'b1, 8'h87, 8'h16}; // CH=6 OP=1
cfg[982] = { 1'b1, 8'h4c, 8'hd}; // CH=3 OP=3
cfg[983] = { 1'b1, 8'h9c, 8'h14}; // CH=3 OP=3
cfg[984] = { 1'b0, 8'h58, 8'h82}; // CH=0 OP=2
cfg[985] = { 1'b0, 8'h84, 8'he3}; // CH=0 OP=1
cfg[986] = { 1'b0, 8'hbf, 8'h27}; // CH=3 OP=3
cfg[987] = { 1'b0, 8'hac, 8'h64}; // CH=0 OP=3
cfg[988] = { 1'b0, 8'h75, 8'h41}; // CH=1 OP=1
cfg[989] = { 1'b1, 8'h58, 8'hf2}; // CH=3 OP=2
cfg[990] = { 1'b0, 8'h3d, 8'h61}; // CH=1 OP=3
cfg[991] = { 1'b1, 8'h53, 8'h82}; // CH=6 OP=0
cfg[992] = { 1'b1, 8'h60, 8'hf1}; // CH=3 OP=0
cfg[993] = { 1'b1, 8'h75, 8'h8}; // CH=4 OP=1
cfg[994] = { 1'b0, 8'hf7, 8'he2}; // CH=3 OP=1
cfg[995] = { 1'b0, 8'hdb, 8'hca}; // CH=3 OP=2
cfg[996] = { 1'b0, 8'haf, 8'he8}; // CH=3 OP=3
cfg[997] = { 1'b1, 8'h5c, 8'h66}; // CH=3 OP=3
cfg[998] = { 1'b1, 8'hd1, 8'ha7}; // CH=4 OP=0
cfg[999] = { 1'b1, 8'hf5, 8'h99}; // CH=4 OP=1
cfg[1000] = { 1'b0, 8'h99, 8'h67}; // CH=1 OP=2
cfg[1001] = { 1'b0, 8'hc4, 8'hba}; // CH=0 OP=1
cfg[1002] = { 1'b1, 8'h3b, 8'h1a}; // CH=6 OP=2
cfg[1003] = { 1'b1, 8'h4f, 8'h8f}; // CH=6 OP=3
cfg[1004] = { 1'b1, 8'hbb, 8'h87}; // CH=6 OP=2
cfg[1005] = { 1'b1, 8'hac, 8'h62}; // CH=3 OP=3
cfg[1006] = { 1'b1, 8'h5b, 8'h64}; // CH=6 OP=2
cfg[1007] = { 1'b0, 8'hb7, 8'hca}; // CH=3 OP=1
cfg[1008] = { 1'b0, 8'h89, 8'h71}; // CH=1 OP=2
cfg[1009] = { 1'b1, 8'hb3, 8'ha}; // CH=6 OP=0
cfg[1010] = { 1'b0, 8'h80, 8'h4}; // CH=0 OP=0
cfg[1011] = { 1'b0, 8'hed, 8'heb}; // CH=1 OP=3
cfg[1012] = { 1'b0, 8'h62, 8'h27}; // CH=2 OP=0
cfg[1013] = { 1'b0, 8'hb9, 8'h76}; // CH=1 OP=2
cfg[1014] = { 1'b1, 8'hda, 8'h32}; // CH=5 OP=2
cfg[1015] = { 1'b1, 8'he3, 8'hde}; // CH=6 OP=0
cfg[1016] = { 1'b1, 8'hd0, 8'h39}; // CH=3 OP=0
cfg[1017] = { 1'b1, 8'hd8, 8'hf1}; // CH=3 OP=2
cfg[1018] = { 1'b0, 8'h71, 8'h7a}; // CH=1 OP=0
cfg[1019] = { 1'b0, 8'hff, 8'h2d}; // CH=3 OP=3
cfg[1020] = { 1'b0, 8'h94, 8'h47}; // CH=0 OP=1
cfg[1021] = { 1'b1, 8'h81, 8'h12}; // CH=4 OP=0
cfg[1022] = { 1'b1, 8'he3, 8'h39}; // CH=6 OP=0
cfg[1023] = { 1'b1, 8'h9c, 8'hb0}; // CH=3 OP=3
cfg[1024] = { 1'b0, 8'h76, 8'he2}; // CH=2 OP=1
cfg[1025] = { 1'b1, 8'h59, 8'hc0}; // CH=4 OP=2
cfg[1026] = { 1'b0, 8'h53, 8'hf9}; // CH=3 OP=0
cfg[1027] = { 1'b0, 8'h59, 8'h1}; // CH=1 OP=2
cfg[1028] = { 1'b0, 8'h69, 8'h72}; // CH=1 OP=2
cfg[1029] = { 1'b1, 8'h7d, 8'h72}; // CH=4 OP=3
cfg[1030] = { 1'b0, 8'hf3, 8'h99}; // CH=3 OP=0
cfg[1031] = { 1'b1, 8'hfd, 8'h92}; // CH=4 OP=3
cfg[1032] = { 1'b1, 8'h84, 8'h75}; // CH=3 OP=1
cfg[1033] = { 1'b1, 8'h77, 8'h11}; // CH=6 OP=1
cfg[1034] = { 1'b1, 8'h37, 8'h4}; // CH=6 OP=1
cfg[1035] = { 1'b1, 8'h30, 8'hc3}; // CH=3 OP=0
cfg[1036] = { 1'b0, 8'h70, 8'h16}; // CH=0 OP=0
cfg[1037] = { 1'b1, 8'hd9, 8'h7e}; // CH=4 OP=2
cfg[1038] = { 1'b1, 8'h57, 8'hf0}; // CH=6 OP=1
cfg[1039] = { 1'b1, 8'h68, 8'h89}; // CH=3 OP=2
cfg[1040] = { 1'b1, 8'hfb, 8'h35}; // CH=6 OP=2
cfg[1041] = { 1'b0, 8'h70, 8'h1a}; // CH=0 OP=0
cfg[1042] = { 1'b0, 8'h82, 8'haf}; // CH=2 OP=0
cfg[1043] = { 1'b1, 8'h74, 8'h26}; // CH=3 OP=1
cfg[1044] = { 1'b1, 8'h37, 8'hea}; // CH=6 OP=1
cfg[1045] = { 1'b1, 8'h4d, 8'hf5}; // CH=4 OP=3
cfg[1046] = { 1'b0, 8'hbd, 8'h1}; // CH=1 OP=3
cfg[1047] = { 1'b0, 8'h97, 8'h7f}; // CH=3 OP=1
cfg[1048] = { 1'b1, 8'hee, 8'h70}; // CH=5 OP=3
cfg[1049] = { 1'b0, 8'h56, 8'hf9}; // CH=2 OP=1
cfg[1050] = { 1'b1, 8'h51, 8'h2e}; // CH=4 OP=0
cfg[1051] = { 1'b1, 8'hc2, 8'h48}; // CH=5 OP=0
cfg[1052] = { 1'b0, 8'h44, 8'hf7}; // CH=0 OP=1
cfg[1053] = { 1'b1, 8'h4d, 8'h1d}; // CH=4 OP=3
cfg[1054] = { 1'b1, 8'h38, 8'h7a}; // CH=3 OP=2
cfg[1055] = { 1'b0, 8'ha0, 8'h8}; // CH=0 OP=0
cfg[1056] = { 1'b0, 8'h5d, 8'h2e}; // CH=1 OP=3
cfg[1057] = { 1'b0, 8'hf4, 8'had}; // CH=0 OP=1
cfg[1058] = { 1'b1, 8'he2, 8'h1d}; // CH=5 OP=0
cfg[1059] = { 1'b0, 8'h39, 8'h17}; // CH=1 OP=2
cfg[1060] = { 1'b1, 8'h8a, 8'h45}; // CH=5 OP=2
cfg[1061] = { 1'b1, 8'h4c, 8'h8e}; // CH=3 OP=3
cfg[1062] = { 1'b1, 8'h90, 8'h85}; // CH=3 OP=0
cfg[1063] = { 1'b0, 8'hde, 8'ha3}; // CH=2 OP=3
cfg[1064] = { 1'b0, 8'h5a, 8'h1d}; // CH=2 OP=2
cfg[1065] = { 1'b1, 8'hfa, 8'h43}; // CH=5 OP=2
cfg[1066] = { 1'b0, 8'h58, 8'h71}; // CH=0 OP=2
cfg[1067] = { 1'b0, 8'h4c, 8'h1e}; // CH=0 OP=3
cfg[1068] = { 1'b0, 8'hf4, 8'h3c}; // CH=0 OP=1
cfg[1069] = { 1'b1, 8'h98, 8'h68}; // CH=3 OP=2
cfg[1070] = { 1'b0, 8'h3f, 8'h34}; // CH=3 OP=3
cfg[1071] = { 1'b1, 8'hcf, 8'hac}; // CH=6 OP=3
cfg[1072] = { 1'b0, 8'had, 8'h4f}; // CH=1 OP=3
cfg[1073] = { 1'b0, 8'hc3, 8'h6c}; // CH=3 OP=0
cfg[1074] = { 1'b0, 8'hc3, 8'h92}; // CH=3 OP=0
cfg[1075] = { 1'b0, 8'h96, 8'h77}; // CH=2 OP=1
cfg[1076] = { 1'b1, 8'hd2, 8'hd6}; // CH=5 OP=0
cfg[1077] = { 1'b0, 8'hfe, 8'hca}; // CH=2 OP=3
cfg[1078] = { 1'b0, 8'hf1, 8'hbd}; // CH=1 OP=0
cfg[1079] = { 1'b0, 8'h30, 8'he4}; // CH=0 OP=0
cfg[1080] = { 1'b0, 8'hff, 8'h90}; // CH=3 OP=3
cfg[1081] = { 1'b0, 8'had, 8'hdf}; // CH=1 OP=3
cfg[1082] = { 1'b0, 8'h70, 8'h4b}; // CH=0 OP=0
cfg[1083] = { 1'b0, 8'h77, 8'hdd}; // CH=3 OP=1
cfg[1084] = { 1'b1, 8'hee, 8'h45}; // CH=5 OP=3
cfg[1085] = { 1'b0, 8'h84, 8'h5c}; // CH=0 OP=1
cfg[1086] = { 1'b0, 8'h56, 8'h32}; // CH=2 OP=1
cfg[1087] = { 1'b0, 8'h7b, 8'hfd}; // CH=3 OP=2
cfg[1088] = { 1'b1, 8'h39, 8'hef}; // CH=4 OP=2
cfg[1089] = { 1'b0, 8'h38, 8'h15}; // CH=0 OP=2
cfg[1090] = { 1'b1, 8'h37, 8'had}; // CH=6 OP=1
cfg[1091] = { 1'b1, 8'he4, 8'h8c}; // CH=3 OP=1
cfg[1092] = { 1'b1, 8'h55, 8'hd7}; // CH=4 OP=1
cfg[1093] = { 1'b0, 8'hcc, 8'hb5}; // CH=0 OP=3
cfg[1094] = { 1'b1, 8'hba, 8'hfa}; // CH=5 OP=2
cfg[1095] = { 1'b0, 8'h3f, 8'h56}; // CH=3 OP=3
cfg[1096] = { 1'b0, 8'h95, 8'h89}; // CH=1 OP=1
cfg[1097] = { 1'b0, 8'h37, 8'h86}; // CH=3 OP=1
cfg[1098] = { 1'b1, 8'h3f, 8'h4a}; // CH=6 OP=3
cfg[1099] = { 1'b0, 8'h77, 8'h67}; // CH=3 OP=1
cfg[1100] = { 1'b0, 8'haf, 8'h14}; // CH=3 OP=3
cfg[1101] = { 1'b1, 8'h93, 8'ha0}; // CH=6 OP=0
cfg[1102] = { 1'b1, 8'he8, 8'h77}; // CH=3 OP=2
cfg[1103] = { 1'b1, 8'hb4, 8'h2c}; // CH=3 OP=1
cfg[1104] = { 1'b0, 8'h6f, 8'h27}; // CH=3 OP=3
cfg[1105] = { 1'b0, 8'hae, 8'h7d}; // CH=2 OP=3
cfg[1106] = { 1'b0, 8'h43, 8'h6}; // CH=3 OP=0
cfg[1107] = { 1'b1, 8'h54, 8'h8c}; // CH=3 OP=1
cfg[1108] = { 1'b0, 8'h9e, 8'h1}; // CH=2 OP=3
cfg[1109] = { 1'b0, 8'h9f, 8'h8c}; // CH=3 OP=3
cfg[1110] = { 1'b0, 8'h4e, 8'h19}; // CH=2 OP=3
cfg[1111] = { 1'b1, 8'he2, 8'hb9}; // CH=5 OP=0
cfg[1112] = { 1'b0, 8'hca, 8'h31}; // CH=2 OP=2
cfg[1113] = { 1'b1, 8'h7f, 8'h5d}; // CH=6 OP=3
cfg[1114] = { 1'b0, 8'hee, 8'h84}; // CH=2 OP=3
cfg[1115] = { 1'b0, 8'h9c, 8'h2}; // CH=0 OP=3
cfg[1116] = { 1'b1, 8'hdf, 8'h8}; // CH=6 OP=3
cfg[1117] = { 1'b0, 8'h34, 8'h95}; // CH=0 OP=1
cfg[1118] = { 1'b0, 8'hd2, 8'h96}; // CH=2 OP=0
cfg[1119] = { 1'b0, 8'hd8, 8'h22}; // CH=0 OP=2
cfg[1120] = { 1'b0, 8'hf1, 8'hee}; // CH=1 OP=0
cfg[1121] = { 1'b0, 8'hab, 8'hb6}; // CH=3 OP=2
cfg[1122] = { 1'b0, 8'hdc, 8'ha8}; // CH=0 OP=3
cfg[1123] = { 1'b1, 8'h39, 8'h32}; // CH=4 OP=2
cfg[1124] = { 1'b0, 8'hbe, 8'hbe}; // CH=2 OP=3
cfg[1125] = { 1'b0, 8'hc0, 8'hd2}; // CH=0 OP=0
cfg[1126] = { 1'b0, 8'hc8, 8'h77}; // CH=0 OP=2
cfg[1127] = { 1'b1, 8'h5d, 8'hcd}; // CH=4 OP=3
cfg[1128] = { 1'b1, 8'hf4, 8'hc}; // CH=3 OP=1
cfg[1129] = { 1'b0, 8'hc8, 8'h72}; // CH=0 OP=2
cfg[1130] = { 1'b0, 8'hb9, 8'h5}; // CH=1 OP=2
cfg[1131] = { 1'b1, 8'h64, 8'hbb}; // CH=3 OP=1
cfg[1132] = { 1'b1, 8'h40, 8'h63}; // CH=3 OP=0
cfg[1133] = { 1'b0, 8'h7a, 8'h95}; // CH=2 OP=2
cfg[1134] = { 1'b0, 8'h38, 8'h53}; // CH=0 OP=2
cfg[1135] = { 1'b0, 8'hf8, 8'h26}; // CH=0 OP=2
cfg[1136] = { 1'b0, 8'hc0, 8'h9d}; // CH=0 OP=0
cfg[1137] = { 1'b0, 8'h77, 8'h6b}; // CH=3 OP=1
cfg[1138] = { 1'b0, 8'he9, 8'hf3}; // CH=1 OP=2
cfg[1139] = { 1'b0, 8'h62, 8'hbb}; // CH=2 OP=0
cfg[1140] = { 1'b1, 8'he8, 8'h75}; // CH=3 OP=2
cfg[1141] = { 1'b1, 8'h4c, 8'h32}; // CH=3 OP=3
cfg[1142] = { 1'b0, 8'he1, 8'h37}; // CH=1 OP=0
cfg[1143] = { 1'b0, 8'h35, 8'hbb}; // CH=1 OP=1
cfg[1144] = { 1'b0, 8'h5b, 8'hae}; // CH=3 OP=2
cfg[1145] = { 1'b0, 8'hf8, 8'haa}; // CH=0 OP=2
cfg[1146] = { 1'b0, 8'h63, 8'h90}; // CH=3 OP=0
cfg[1147] = { 1'b0, 8'hda, 8'h94}; // CH=2 OP=2
cfg[1148] = { 1'b0, 8'hc4, 8'h87}; // CH=0 OP=1
cfg[1149] = { 1'b1, 8'hb8, 8'h43}; // CH=3 OP=2
cfg[1150] = { 1'b1, 8'h91, 8'hf3}; // CH=4 OP=0
cfg[1151] = { 1'b1, 8'hab, 8'h3f}; // CH=6 OP=2
cfg[1152] = { 1'b0, 8'h3f, 8'h20}; // CH=3 OP=3
cfg[1153] = { 1'b0, 8'hb0, 8'h55}; // CH=0 OP=0
cfg[1154] = { 1'b1, 8'ha9, 8'hd2}; // CH=4 OP=2
cfg[1155] = { 1'b0, 8'hf6, 8'h63}; // CH=2 OP=1
cfg[1156] = { 1'b1, 8'hab, 8'he7}; // CH=6 OP=2
cfg[1157] = { 1'b0, 8'h88, 8'hab}; // CH=0 OP=2
cfg[1158] = { 1'b1, 8'h92, 8'hd1}; // CH=5 OP=0
cfg[1159] = { 1'b1, 8'h85, 8'h26}; // CH=4 OP=1
cfg[1160] = { 1'b1, 8'hc4, 8'had}; // CH=3 OP=1
cfg[1161] = { 1'b0, 8'he5, 8'h6c}; // CH=1 OP=1
cfg[1162] = { 1'b0, 8'h3a, 8'he6}; // CH=2 OP=2
cfg[1163] = { 1'b1, 8'heb, 8'he}; // CH=6 OP=2
cfg[1164] = { 1'b1, 8'h94, 8'he0}; // CH=3 OP=1
cfg[1165] = { 1'b1, 8'ha0, 8'h43}; // CH=3 OP=0
cfg[1166] = { 1'b1, 8'h87, 8'h3a}; // CH=6 OP=1
cfg[1167] = { 1'b0, 8'h32, 8'hb9}; // CH=2 OP=0
cfg[1168] = { 1'b0, 8'he1, 8'h7a}; // CH=1 OP=0
cfg[1169] = { 1'b0, 8'h66, 8'h29}; // CH=2 OP=1
cfg[1170] = { 1'b1, 8'hb5, 8'hd7}; // CH=4 OP=1
cfg[1171] = { 1'b1, 8'hab, 8'h10}; // CH=6 OP=2
cfg[1172] = { 1'b1, 8'had, 8'h4a}; // CH=4 OP=3
cfg[1173] = { 1'b1, 8'h7e, 8'h35}; // CH=5 OP=3
cfg[1174] = { 1'b1, 8'ha3, 8'hc9}; // CH=6 OP=0
cfg[1175] = { 1'b1, 8'hbe, 8'h6a}; // CH=5 OP=3
cfg[1176] = { 1'b1, 8'h85, 8'hf1}; // CH=4 OP=1
cfg[1177] = { 1'b0, 8'hd3, 8'h24}; // CH=3 OP=0
cfg[1178] = { 1'b1, 8'hb4, 8'h27}; // CH=3 OP=1
cfg[1179] = { 1'b1, 8'hbc, 8'h51}; // CH=3 OP=3
cfg[1180] = { 1'b0, 8'h71, 8'h46}; // CH=1 OP=0
cfg[1181] = { 1'b1, 8'h94, 8'h56}; // CH=3 OP=1
cfg[1182] = { 1'b0, 8'hcb, 8'hca}; // CH=3 OP=2
cfg[1183] = { 1'b0, 8'he2, 8'h48}; // CH=2 OP=0
cfg[1184] = { 1'b1, 8'h3d, 8'heb}; // CH=4 OP=3
cfg[1185] = { 1'b1, 8'hd3, 8'ha9}; // CH=6 OP=0
cfg[1186] = { 1'b1, 8'hea, 8'h2e}; // CH=5 OP=2
cfg[1187] = { 1'b0, 8'ha7, 8'hb6}; // CH=3 OP=1
cfg[1188] = { 1'b1, 8'h63, 8'hd1}; // CH=6 OP=0
cfg[1189] = { 1'b1, 8'hd5, 8'h17}; // CH=4 OP=1
cfg[1190] = { 1'b0, 8'hf2, 8'h6d}; // CH=2 OP=0
cfg[1191] = { 1'b0, 8'hbc, 8'he}; // CH=0 OP=3
cfg[1192] = { 1'b1, 8'h6c, 8'he4}; // CH=3 OP=3
cfg[1193] = { 1'b1, 8'ha9, 8'hef}; // CH=4 OP=2
cfg[1194] = { 1'b1, 8'h7c, 8'h98}; // CH=3 OP=3
cfg[1195] = { 1'b0, 8'h9e, 8'hc7}; // CH=2 OP=3
cfg[1196] = { 1'b1, 8'h88, 8'hc9}; // CH=3 OP=2
cfg[1197] = { 1'b1, 8'h30, 8'h7f}; // CH=3 OP=0
cfg[1198] = { 1'b1, 8'h93, 8'h51}; // CH=6 OP=0
cfg[1199] = { 1'b0, 8'h68, 8'h68}; // CH=0 OP=2
cfg[1200] = { 1'b1, 8'h5a, 8'hd6}; // CH=5 OP=2
cfg[1201] = { 1'b1, 8'hb7, 8'he4}; // CH=6 OP=1
cfg[1202] = { 1'b0, 8'h4b, 8'h1a}; // CH=3 OP=2
cfg[1203] = { 1'b1, 8'hd8, 8'hcc}; // CH=3 OP=2
cfg[1204] = { 1'b0, 8'h60, 8'h49}; // CH=0 OP=0
cfg[1205] = { 1'b1, 8'h32, 8'he7}; // CH=5 OP=0
cfg[1206] = { 1'b1, 8'hb1, 8'hf5}; // CH=4 OP=0
cfg[1207] = { 1'b1, 8'h33, 8'h7a}; // CH=6 OP=0
cfg[1208] = { 1'b0, 8'h9b, 8'h6b}; // CH=3 OP=2
cfg[1209] = { 1'b1, 8'hf6, 8'h41}; // CH=5 OP=1
cfg[1210] = { 1'b1, 8'hed, 8'h25}; // CH=4 OP=3
cfg[1211] = { 1'b1, 8'h38, 8'h35}; // CH=3 OP=2
cfg[1212] = { 1'b0, 8'hd2, 8'h1}; // CH=2 OP=0
cfg[1213] = { 1'b0, 8'h3b, 8'h71}; // CH=3 OP=2
cfg[1214] = { 1'b1, 8'h6d, 8'h79}; // CH=4 OP=3
cfg[1215] = { 1'b1, 8'h40, 8'h6e}; // CH=3 OP=0
cfg[1216] = { 1'b0, 8'h73, 8'h21}; // CH=3 OP=0
cfg[1217] = { 1'b0, 8'hd4, 8'h8c}; // CH=0 OP=1
cfg[1218] = { 1'b1, 8'hf2, 8'h5}; // CH=5 OP=0
cfg[1219] = { 1'b1, 8'hdf, 8'h41}; // CH=6 OP=3
cfg[1220] = { 1'b0, 8'h69, 8'h76}; // CH=1 OP=2
cfg[1221] = { 1'b1, 8'h3b, 8'h29}; // CH=6 OP=2
cfg[1222] = { 1'b0, 8'h77, 8'h9a}; // CH=3 OP=1
cfg[1223] = { 1'b1, 8'he4, 8'h13}; // CH=3 OP=1
cfg[1224] = { 1'b0, 8'hd5, 8'h81}; // CH=1 OP=1
cfg[1225] = { 1'b1, 8'h48, 8'h25}; // CH=3 OP=2
cfg[1226] = { 1'b0, 8'h57, 8'hb1}; // CH=3 OP=1
cfg[1227] = { 1'b0, 8'h5c, 8'h7f}; // CH=0 OP=3
cfg[1228] = { 1'b1, 8'h6e, 8'h71}; // CH=5 OP=3
cfg[1229] = { 1'b0, 8'ha6, 8'h51}; // CH=2 OP=1
cfg[1230] = { 1'b0, 8'h41, 8'h69}; // CH=1 OP=0
cfg[1231] = { 1'b0, 8'hc2, 8'h4b}; // CH=2 OP=0
cfg[1232] = { 1'b1, 8'ha6, 8'h40}; // CH=5 OP=1
cfg[1233] = { 1'b1, 8'haa, 8'hc1}; // CH=5 OP=2
cfg[1234] = { 1'b0, 8'hcf, 8'h2b}; // CH=3 OP=3
cfg[1235] = { 1'b1, 8'h80, 8'h3b}; // CH=3 OP=0
cfg[1236] = { 1'b0, 8'hff, 8'h1f}; // CH=3 OP=3
cfg[1237] = { 1'b1, 8'h71, 8'h32}; // CH=4 OP=0
cfg[1238] = { 1'b1, 8'hc2, 8'h86}; // CH=5 OP=0
cfg[1239] = { 1'b1, 8'h81, 8'h50}; // CH=4 OP=0
cfg[1240] = { 1'b1, 8'hcc, 8'hbd}; // CH=3 OP=3
cfg[1241] = { 1'b1, 8'h8e, 8'he9}; // CH=5 OP=3
cfg[1242] = { 1'b0, 8'h34, 8'h29}; // CH=0 OP=1
cfg[1243] = { 1'b1, 8'hde, 8'heb}; // CH=5 OP=3
cfg[1244] = { 1'b0, 8'had, 8'h16}; // CH=1 OP=3
cfg[1245] = { 1'b1, 8'h70, 8'h51}; // CH=3 OP=0
cfg[1246] = { 1'b1, 8'ha2, 8'h7e}; // CH=5 OP=0
cfg[1247] = { 1'b0, 8'h60, 8'h49}; // CH=0 OP=0
cfg[1248] = { 1'b1, 8'h8b, 8'h78}; // CH=6 OP=2
cfg[1249] = { 1'b0, 8'h48, 8'h9}; // CH=0 OP=2
cfg[1250] = { 1'b0, 8'h32, 8'h9e}; // CH=2 OP=0
cfg[1251] = { 1'b0, 8'h5b, 8'h2a}; // CH=3 OP=2
cfg[1252] = { 1'b0, 8'h46, 8'h42}; // CH=2 OP=1
cfg[1253] = { 1'b1, 8'h5c, 8'hba}; // CH=3 OP=3
cfg[1254] = { 1'b0, 8'had, 8'hdb}; // CH=1 OP=3
cfg[1255] = { 1'b0, 8'hb2, 8'hfc}; // CH=2 OP=0
cfg[1256] = { 1'b1, 8'h50, 8'hbf}; // CH=3 OP=0
cfg[1257] = { 1'b0, 8'hb1, 8'he7}; // CH=1 OP=0
cfg[1258] = { 1'b1, 8'h3c, 8'h5f}; // CH=3 OP=3
cfg[1259] = { 1'b1, 8'h85, 8'h69}; // CH=4 OP=1
cfg[1260] = { 1'b1, 8'hb7, 8'h7}; // CH=6 OP=1
cfg[1261] = { 1'b1, 8'h74, 8'h32}; // CH=3 OP=1
cfg[1262] = { 1'b1, 8'hb5, 8'hcd}; // CH=4 OP=1
cfg[1263] = { 1'b1, 8'h63, 8'h9}; // CH=6 OP=0
cfg[1264] = { 1'b0, 8'h80, 8'h5}; // CH=0 OP=0
cfg[1265] = { 1'b0, 8'h40, 8'h80}; // CH=0 OP=0
cfg[1266] = { 1'b0, 8'h5b, 8'h45}; // CH=3 OP=2
cfg[1267] = { 1'b0, 8'h98, 8'h87}; // CH=0 OP=2
cfg[1268] = { 1'b0, 8'h43, 8'hf0}; // CH=3 OP=0
cfg[1269] = { 1'b1, 8'h9d, 8'hd4}; // CH=4 OP=3
cfg[1270] = { 1'b1, 8'hc1, 8'he6}; // CH=4 OP=0
cfg[1271] = { 1'b1, 8'h8e, 8'h3f}; // CH=5 OP=3
cfg[1272] = { 1'b1, 8'hb1, 8'hf5}; // CH=4 OP=0
cfg[1273] = { 1'b0, 8'h59, 8'h58}; // CH=1 OP=2
cfg[1274] = { 1'b0, 8'hb3, 8'hd8}; // CH=3 OP=0
cfg[1275] = { 1'b0, 8'h5e, 8'h18}; // CH=2 OP=3
cfg[1276] = { 1'b1, 8'hb9, 8'h40}; // CH=4 OP=2
cfg[1277] = { 1'b0, 8'h51, 8'hc7}; // CH=1 OP=0
cfg[1278] = { 1'b0, 8'h6e, 8'hb7}; // CH=2 OP=3
cfg[1279] = { 1'b1, 8'h42, 8'hae}; // CH=5 OP=0
cfg[1280] = { 1'b0, 8'h85, 8'hd8}; // CH=1 OP=1
cfg[1281] = { 1'b1, 8'h41, 8'h68}; // CH=4 OP=0
cfg[1282] = { 1'b1, 8'hb5, 8'hc5}; // CH=4 OP=1
cfg[1283] = { 1'b0, 8'h8e, 8'hef}; // CH=2 OP=3
cfg[1284] = { 1'b0, 8'ha6, 8'h4a}; // CH=2 OP=1
cfg[1285] = { 1'b0, 8'he6, 8'he9}; // CH=2 OP=1
cfg[1286] = { 1'b1, 8'had, 8'h4d}; // CH=4 OP=3
cfg[1287] = { 1'b1, 8'h64, 8'h31}; // CH=3 OP=1
cfg[1288] = { 1'b1, 8'hec, 8'h59}; // CH=3 OP=3
cfg[1289] = { 1'b1, 8'ha3, 8'heb}; // CH=6 OP=0
cfg[1290] = { 1'b0, 8'hb6, 8'h7d}; // CH=2 OP=1
cfg[1291] = { 1'b1, 8'h7b, 8'hdb}; // CH=6 OP=2
cfg[1292] = { 1'b1, 8'h9a, 8'h90}; // CH=5 OP=2
cfg[1293] = { 1'b0, 8'h6c, 8'h1e}; // CH=0 OP=3
cfg[1294] = { 1'b0, 8'h9c, 8'hc5}; // CH=0 OP=3
cfg[1295] = { 1'b0, 8'h85, 8'hab}; // CH=1 OP=1
cfg[1296] = { 1'b1, 8'hc0, 8'h59}; // CH=3 OP=0
cfg[1297] = { 1'b1, 8'h6a, 8'hbd}; // CH=5 OP=2
cfg[1298] = { 1'b0, 8'h56, 8'hd0}; // CH=2 OP=1
cfg[1299] = { 1'b1, 8'h6b, 8'hbb}; // CH=6 OP=2
cfg[1300] = { 1'b0, 8'he8, 8'h1c}; // CH=0 OP=2
cfg[1301] = { 1'b1, 8'hc3, 8'hbd}; // CH=6 OP=0
cfg[1302] = { 1'b0, 8'h54, 8'h74}; // CH=0 OP=1
cfg[1303] = { 1'b0, 8'h72, 8'h1b}; // CH=2 OP=0
cfg[1304] = { 1'b0, 8'h37, 8'hb}; // CH=3 OP=1
cfg[1305] = { 1'b0, 8'he3, 8'he5}; // CH=3 OP=0
cfg[1306] = { 1'b0, 8'h3c, 8'hd}; // CH=0 OP=3
cfg[1307] = { 1'b0, 8'hf9, 8'h66}; // CH=1 OP=2
cfg[1308] = { 1'b0, 8'hca, 8'h18}; // CH=2 OP=2
cfg[1309] = { 1'b0, 8'h85, 8'he7}; // CH=1 OP=1
cfg[1310] = { 1'b1, 8'ha1, 8'h5a}; // CH=4 OP=0
cfg[1311] = { 1'b0, 8'h5f, 8'h83}; // CH=3 OP=3
cfg[1312] = { 1'b1, 8'hd3, 8'h27}; // CH=6 OP=0
cfg[1313] = { 1'b1, 8'hee, 8'h66}; // CH=5 OP=3
cfg[1314] = { 1'b0, 8'hfa, 8'h10}; // CH=2 OP=2
cfg[1315] = { 1'b1, 8'hdf, 8'h57}; // CH=6 OP=3
cfg[1316] = { 1'b0, 8'hec, 8'h23}; // CH=0 OP=3
cfg[1317] = { 1'b0, 8'h52, 8'haf}; // CH=2 OP=0
cfg[1318] = { 1'b0, 8'h6a, 8'ha6}; // CH=2 OP=2
cfg[1319] = { 1'b0, 8'h52, 8'hf2}; // CH=2 OP=0
cfg[1320] = { 1'b1, 8'hac, 8'haa}; // CH=3 OP=3
cfg[1321] = { 1'b1, 8'hca, 8'h4a}; // CH=5 OP=2
cfg[1322] = { 1'b1, 8'h9d, 8'h56}; // CH=4 OP=3
cfg[1323] = { 1'b1, 8'h8c, 8'hbc}; // CH=3 OP=3
cfg[1324] = { 1'b1, 8'h86, 8'hcd}; // CH=5 OP=1
cfg[1325] = { 1'b0, 8'h65, 8'h24}; // CH=1 OP=1
cfg[1326] = { 1'b1, 8'h52, 8'h47}; // CH=5 OP=0
cfg[1327] = { 1'b1, 8'ha4, 8'hf6}; // CH=3 OP=1
cfg[1328] = { 1'b1, 8'h73, 8'h9c}; // CH=6 OP=0
cfg[1329] = { 1'b1, 8'h3d, 8'h61}; // CH=4 OP=3
cfg[1330] = { 1'b1, 8'ha8, 8'hd}; // CH=3 OP=2
cfg[1331] = { 1'b1, 8'h72, 8'h3c}; // CH=5 OP=0
cfg[1332] = { 1'b0, 8'h95, 8'h92}; // CH=1 OP=1
cfg[1333] = { 1'b1, 8'h40, 8'h9b}; // CH=3 OP=0
cfg[1334] = { 1'b1, 8'h87, 8'h4a}; // CH=6 OP=1
cfg[1335] = { 1'b1, 8'h7d, 8'hff}; // CH=4 OP=3
cfg[1336] = { 1'b1, 8'h8c, 8'h2f}; // CH=3 OP=3
cfg[1337] = { 1'b0, 8'hed, 8'ha9}; // CH=1 OP=3
cfg[1338] = { 1'b1, 8'hfa, 8'he2}; // CH=5 OP=2
cfg[1339] = { 1'b1, 8'h36, 8'h65}; // CH=5 OP=1
cfg[1340] = { 1'b1, 8'hc9, 8'h95}; // CH=4 OP=2
cfg[1341] = { 1'b1, 8'ha4, 8'h2b}; // CH=3 OP=1
cfg[1342] = { 1'b1, 8'hc6, 8'h34}; // CH=5 OP=1
cfg[1343] = { 1'b0, 8'h4d, 8'h74}; // CH=1 OP=3
cfg[1344] = { 1'b0, 8'hae, 8'hfb}; // CH=2 OP=3
cfg[1345] = { 1'b0, 8'hdd, 8'ha3}; // CH=1 OP=3
cfg[1346] = { 1'b0, 8'h7f, 8'h30}; // CH=3 OP=3
cfg[1347] = { 1'b1, 8'h5f, 8'h1d}; // CH=6 OP=3
cfg[1348] = { 1'b1, 8'he6, 8'h18}; // CH=5 OP=1
cfg[1349] = { 1'b0, 8'he0, 8'h4e}; // CH=0 OP=0
cfg[1350] = { 1'b0, 8'he9, 8'h17}; // CH=1 OP=2
cfg[1351] = { 1'b1, 8'h8d, 8'h2f}; // CH=4 OP=3
cfg[1352] = { 1'b0, 8'h53, 8'h63}; // CH=3 OP=0
cfg[1353] = { 1'b1, 8'ha0, 8'hd7}; // CH=3 OP=0
cfg[1354] = { 1'b1, 8'hc6, 8'hd2}; // CH=5 OP=1
cfg[1355] = { 1'b1, 8'h6a, 8'h4b}; // CH=5 OP=2
cfg[1356] = { 1'b0, 8'h9a, 8'hdd}; // CH=2 OP=2
cfg[1357] = { 1'b0, 8'hb7, 8'h19}; // CH=3 OP=1
cfg[1358] = { 1'b1, 8'hcf, 8'h36}; // CH=6 OP=3
cfg[1359] = { 1'b1, 8'hd5, 8'hb9}; // CH=4 OP=1
cfg[1360] = { 1'b1, 8'hbe, 8'h35}; // CH=5 OP=3
cfg[1361] = { 1'b0, 8'h4c, 8'h65}; // CH=0 OP=3
cfg[1362] = { 1'b0, 8'h9f, 8'hc8}; // CH=3 OP=3
cfg[1363] = { 1'b1, 8'h40, 8'ha0}; // CH=3 OP=0
cfg[1364] = { 1'b1, 8'h96, 8'h72}; // CH=5 OP=1
cfg[1365] = { 1'b1, 8'hc7, 8'h70}; // CH=6 OP=1
cfg[1366] = { 1'b1, 8'h77, 8'ha}; // CH=6 OP=1
cfg[1367] = { 1'b0, 8'h86, 8'hc2}; // CH=2 OP=1
cfg[1368] = { 1'b0, 8'h7b, 8'h91}; // CH=3 OP=2
cfg[1369] = { 1'b1, 8'h51, 8'haf}; // CH=4 OP=0
cfg[1370] = { 1'b0, 8'h88, 8'he5}; // CH=0 OP=2
cfg[1371] = { 1'b0, 8'hfb, 8'h5b}; // CH=3 OP=2
cfg[1372] = { 1'b0, 8'h3b, 8'hb2}; // CH=3 OP=2
cfg[1373] = { 1'b1, 8'h41, 8'h25}; // CH=4 OP=0
cfg[1374] = { 1'b0, 8'hb2, 8'he2}; // CH=2 OP=0
cfg[1375] = { 1'b1, 8'hbc, 8'h7d}; // CH=3 OP=3
cfg[1376] = { 1'b0, 8'h7e, 8'h31}; // CH=2 OP=3
cfg[1377] = { 1'b0, 8'he5, 8'h1c}; // CH=1 OP=1
cfg[1378] = { 1'b1, 8'h36, 8'hbf}; // CH=5 OP=1
cfg[1379] = { 1'b0, 8'h46, 8'ha4}; // CH=2 OP=1
cfg[1380] = { 1'b0, 8'ha1, 8'hee}; // CH=1 OP=0
cfg[1381] = { 1'b1, 8'h9c, 8'h1}; // CH=3 OP=3
cfg[1382] = { 1'b0, 8'hd7, 8'hb3}; // CH=3 OP=1
cfg[1383] = { 1'b1, 8'h6d, 8'hd8}; // CH=4 OP=3
cfg[1384] = { 1'b1, 8'hda, 8'hcb}; // CH=5 OP=2
cfg[1385] = { 1'b0, 8'hbe, 8'h87}; // CH=2 OP=3
cfg[1386] = { 1'b0, 8'h86, 8'h6}; // CH=2 OP=1
cfg[1387] = { 1'b0, 8'h45, 8'he}; // CH=1 OP=1
cfg[1388] = { 1'b1, 8'h79, 8'h44}; // CH=4 OP=2
cfg[1389] = { 1'b0, 8'h36, 8'h8a}; // CH=2 OP=1
cfg[1390] = { 1'b0, 8'h69, 8'h2c}; // CH=1 OP=2
cfg[1391] = { 1'b0, 8'ha0, 8'hd9}; // CH=0 OP=0
cfg[1392] = { 1'b1, 8'hb9, 8'hf5}; // CH=4 OP=2
cfg[1393] = { 1'b0, 8'h84, 8'hb0}; // CH=0 OP=1
cfg[1394] = { 1'b1, 8'ha7, 8'he9}; // CH=6 OP=1
cfg[1395] = { 1'b1, 8'hd0, 8'h11}; // CH=3 OP=0
cfg[1396] = { 1'b1, 8'hde, 8'h27}; // CH=5 OP=3
cfg[1397] = { 1'b0, 8'h98, 8'hfd}; // CH=0 OP=2
cfg[1398] = { 1'b1, 8'hce, 8'had}; // CH=5 OP=3
cfg[1399] = { 1'b1, 8'hef, 8'hd9}; // CH=6 OP=3
cfg[1400] = { 1'b1, 8'hc9, 8'ha1}; // CH=4 OP=2
cfg[1401] = { 1'b0, 8'h6a, 8'h41}; // CH=2 OP=2
cfg[1402] = { 1'b1, 8'h78, 8'hfa}; // CH=3 OP=2
cfg[1403] = { 1'b0, 8'h61, 8'h7e}; // CH=1 OP=0
cfg[1404] = { 1'b1, 8'h48, 8'h8a}; // CH=3 OP=2
cfg[1405] = { 1'b1, 8'hc3, 8'hd9}; // CH=6 OP=0
cfg[1406] = { 1'b1, 8'hc0, 8'h3f}; // CH=3 OP=0
cfg[1407] = { 1'b1, 8'h37, 8'hd7}; // CH=6 OP=1
cfg[1408] = { 1'b0, 8'h5f, 8'ha5}; // CH=3 OP=3
cfg[1409] = { 1'b1, 8'h5e, 8'h5f}; // CH=5 OP=3
cfg[1410] = { 1'b1, 8'hc8, 8'h42}; // CH=3 OP=2
cfg[1411] = { 1'b1, 8'h40, 8'h3d}; // CH=3 OP=0
cfg[1412] = { 1'b1, 8'ha2, 8'hbb}; // CH=5 OP=0
cfg[1413] = { 1'b0, 8'hab, 8'h45}; // CH=3 OP=2
cfg[1414] = { 1'b0, 8'h84, 8'he1}; // CH=0 OP=1
cfg[1415] = { 1'b1, 8'h3b, 8'ha4}; // CH=6 OP=2
cfg[1416] = { 1'b0, 8'ha2, 8'h64}; // CH=2 OP=0
cfg[1417] = { 1'b1, 8'h47, 8'h9b}; // CH=6 OP=1
cfg[1418] = { 1'b1, 8'hdc, 8'hfa}; // CH=3 OP=3
cfg[1419] = { 1'b1, 8'h3a, 8'hfb}; // CH=5 OP=2
cfg[1420] = { 1'b0, 8'hf7, 8'h3e}; // CH=3 OP=1
cfg[1421] = { 1'b1, 8'h36, 8'h43}; // CH=5 OP=1
cfg[1422] = { 1'b1, 8'h7c, 8'h46}; // CH=3 OP=3
cfg[1423] = { 1'b0, 8'h5d, 8'hb0}; // CH=1 OP=3
cfg[1424] = { 1'b0, 8'h4f, 8'h3b}; // CH=3 OP=3
cfg[1425] = { 1'b0, 8'h63, 8'h65}; // CH=3 OP=0
cfg[1426] = { 1'b0, 8'hfe, 8'h0}; // CH=2 OP=3
cfg[1427] = { 1'b1, 8'hf9, 8'hb1}; // CH=4 OP=2
cfg[1428] = { 1'b0, 8'hf4, 8'hc2}; // CH=0 OP=1
cfg[1429] = { 1'b0, 8'h32, 8'h99}; // CH=2 OP=0
cfg[1430] = { 1'b1, 8'had, 8'h90}; // CH=4 OP=3
cfg[1431] = { 1'b0, 8'he4, 8'hb5}; // CH=0 OP=1
cfg[1432] = { 1'b1, 8'h60, 8'hfb}; // CH=3 OP=0
cfg[1433] = { 1'b1, 8'hbd, 8'hac}; // CH=4 OP=3
cfg[1434] = { 1'b1, 8'hbe, 8'he7}; // CH=5 OP=3
cfg[1435] = { 1'b0, 8'h87, 8'hed}; // CH=3 OP=1
cfg[1436] = { 1'b1, 8'h86, 8'h23}; // CH=5 OP=1
cfg[1437] = { 1'b1, 8'h7f, 8'hd4}; // CH=6 OP=3
cfg[1438] = { 1'b1, 8'h73, 8'h97}; // CH=6 OP=0
cfg[1439] = { 1'b1, 8'ha6, 8'h30}; // CH=5 OP=1
cfg[1440] = { 1'b0, 8'h53, 8'hc0}; // CH=3 OP=0
cfg[1441] = { 1'b0, 8'h37, 8'h75}; // CH=3 OP=1
cfg[1442] = { 1'b1, 8'h97, 8'h71}; // CH=6 OP=1
cfg[1443] = { 1'b0, 8'h54, 8'h1d}; // CH=0 OP=1
cfg[1444] = { 1'b1, 8'h97, 8'h4}; // CH=6 OP=1
cfg[1445] = { 1'b0, 8'h87, 8'h35}; // CH=3 OP=1
cfg[1446] = { 1'b0, 8'h5d, 8'ha5}; // CH=1 OP=3
cfg[1447] = { 1'b0, 8'hb5, 8'h97}; // CH=1 OP=1
cfg[1448] = { 1'b0, 8'hb4, 8'h3d}; // CH=0 OP=1
cfg[1449] = { 1'b1, 8'hc8, 8'hc2}; // CH=3 OP=2
cfg[1450] = { 1'b1, 8'h60, 8'h9b}; // CH=3 OP=0
cfg[1451] = { 1'b0, 8'hb4, 8'hb8}; // CH=0 OP=1
cfg[1452] = { 1'b1, 8'hc7, 8'hbc}; // CH=6 OP=1
cfg[1453] = { 1'b1, 8'hfc, 8'hae}; // CH=3 OP=3
cfg[1454] = { 1'b0, 8'h55, 8'h36}; // CH=1 OP=1
cfg[1455] = { 1'b1, 8'h82, 8'h42}; // CH=5 OP=0
cfg[1456] = { 1'b1, 8'h46, 8'ha0}; // CH=5 OP=1
cfg[1457] = { 1'b0, 8'h3a, 8'h55}; // CH=2 OP=2
cfg[1458] = { 1'b0, 8'hee, 8'h6a}; // CH=2 OP=3
cfg[1459] = { 1'b1, 8'h5f, 8'h2c}; // CH=6 OP=3
cfg[1460] = { 1'b0, 8'hbf, 8'hb3}; // CH=3 OP=3
cfg[1461] = { 1'b0, 8'h74, 8'h6b}; // CH=0 OP=1
cfg[1462] = { 1'b1, 8'h3b, 8'h28}; // CH=6 OP=2
cfg[1463] = { 1'b0, 8'h37, 8'hd6}; // CH=3 OP=1
cfg[1464] = { 1'b0, 8'h8c, 8'hc}; // CH=0 OP=3
cfg[1465] = { 1'b1, 8'haa, 8'h4f}; // CH=5 OP=2
cfg[1466] = { 1'b1, 8'h73, 8'h54}; // CH=6 OP=0
cfg[1467] = { 1'b0, 8'h79, 8'h8e}; // CH=1 OP=2
cfg[1468] = { 1'b0, 8'hdb, 8'h7d}; // CH=3 OP=2
cfg[1469] = { 1'b1, 8'ha7, 8'h6f}; // CH=6 OP=1
cfg[1470] = { 1'b1, 8'hb1, 8'h2f}; // CH=4 OP=0
cfg[1471] = { 1'b0, 8'h6c, 8'ha3}; // CH=0 OP=3
cfg[1472] = { 1'b0, 8'h71, 8'hde}; // CH=1 OP=0
cfg[1473] = { 1'b1, 8'hdd, 8'h15}; // CH=4 OP=3
cfg[1474] = { 1'b1, 8'h57, 8'ha2}; // CH=6 OP=1
cfg[1475] = { 1'b0, 8'hfd, 8'hb0}; // CH=1 OP=3
cfg[1476] = { 1'b1, 8'h41, 8'h74}; // CH=4 OP=0
cfg[1477] = { 1'b1, 8'hf0, 8'hed}; // CH=3 OP=0
cfg[1478] = { 1'b0, 8'hcb, 8'hfd}; // CH=3 OP=2
cfg[1479] = { 1'b0, 8'h72, 8'h6d}; // CH=2 OP=0
cfg[1480] = { 1'b1, 8'ha3, 8'h9c}; // CH=6 OP=0
cfg[1481] = { 1'b1, 8'h80, 8'h8f}; // CH=3 OP=0
cfg[1482] = { 1'b1, 8'h33, 8'h0}; // CH=6 OP=0
cfg[1483] = { 1'b0, 8'hf2, 8'hde}; // CH=2 OP=0
cfg[1484] = { 1'b0, 8'h85, 8'h35}; // CH=1 OP=1
cfg[1485] = { 1'b0, 8'h8a, 8'hfe}; // CH=2 OP=2
cfg[1486] = { 1'b1, 8'h98, 8'h40}; // CH=3 OP=2
cfg[1487] = { 1'b0, 8'h96, 8'h2e}; // CH=2 OP=1
cfg[1488] = { 1'b1, 8'h6d, 8'hd4}; // CH=4 OP=3
cfg[1489] = { 1'b1, 8'h90, 8'h9f}; // CH=3 OP=0
cfg[1490] = { 1'b0, 8'he6, 8'hde}; // CH=2 OP=1
cfg[1491] = { 1'b1, 8'hfe, 8'h20}; // CH=5 OP=3
cfg[1492] = { 1'b0, 8'h33, 8'h2}; // CH=3 OP=0
cfg[1493] = { 1'b1, 8'h69, 8'h87}; // CH=4 OP=2
cfg[1494] = { 1'b1, 8'h4b, 8'h11}; // CH=6 OP=2
cfg[1495] = { 1'b0, 8'h7b, 8'had}; // CH=3 OP=2
cfg[1496] = { 1'b0, 8'h76, 8'h43}; // CH=2 OP=1
cfg[1497] = { 1'b0, 8'he3, 8'h46}; // CH=3 OP=0
cfg[1498] = { 1'b1, 8'h73, 8'he5}; // CH=6 OP=0
cfg[1499] = { 1'b0, 8'h93, 8'hc3}; // CH=3 OP=0
cfg[1500] = { 1'b0, 8'hb3, 8'hbe}; // CH=3 OP=0
cfg[1501] = { 1'b0, 8'hb1, 8'heb}; // CH=1 OP=0
cfg[1502] = { 1'b0, 8'he4, 8'hed}; // CH=0 OP=1
cfg[1503] = { 1'b1, 8'h4d, 8'h74}; // CH=4 OP=3
cfg[1504] = { 1'b0, 8'h62, 8'h85}; // CH=2 OP=0
cfg[1505] = { 1'b0, 8'h45, 8'hb4}; // CH=1 OP=1
cfg[1506] = { 1'b0, 8'hbc, 8'h52}; // CH=0 OP=3
cfg[1507] = { 1'b1, 8'h9f, 8'h98}; // CH=6 OP=3
cfg[1508] = { 1'b0, 8'h8e, 8'h7d}; // CH=2 OP=3
cfg[1509] = { 1'b0, 8'hcf, 8'ha6}; // CH=3 OP=3
cfg[1510] = { 1'b0, 8'he9, 8'h59}; // CH=1 OP=2
cfg[1511] = { 1'b0, 8'hd7, 8'h8f}; // CH=3 OP=1
cfg[1512] = { 1'b0, 8'h4b, 8'h2}; // CH=3 OP=2
cfg[1513] = { 1'b1, 8'hd1, 8'h80}; // CH=4 OP=0
cfg[1514] = { 1'b1, 8'h85, 8'h4a}; // CH=4 OP=1
cfg[1515] = { 1'b0, 8'h95, 8'h90}; // CH=1 OP=1
cfg[1516] = { 1'b0, 8'hd6, 8'h4c}; // CH=2 OP=1
cfg[1517] = { 1'b0, 8'hfe, 8'heb}; // CH=2 OP=3
cfg[1518] = { 1'b1, 8'ha4, 8'h53}; // CH=3 OP=1
cfg[1519] = { 1'b0, 8'hfd, 8'h51}; // CH=1 OP=3
cfg[1520] = { 1'b1, 8'hf5, 8'h3b}; // CH=4 OP=1
cfg[1521] = { 1'b0, 8'h31, 8'h5d}; // CH=1 OP=0
cfg[1522] = { 1'b1, 8'hce, 8'h2e}; // CH=5 OP=3
cfg[1523] = { 1'b1, 8'h7b, 8'hb3}; // CH=6 OP=2
cfg[1524] = { 1'b1, 8'h79, 8'h49}; // CH=4 OP=2
cfg[1525] = { 1'b1, 8'hb5, 8'h1f}; // CH=4 OP=1
cfg[1526] = { 1'b0, 8'hb3, 8'h23}; // CH=3 OP=0
cfg[1527] = { 1'b0, 8'h58, 8'h77}; // CH=0 OP=2
cfg[1528] = { 1'b0, 8'h55, 8'hc8}; // CH=1 OP=1
cfg[1529] = { 1'b0, 8'h5d, 8'h3}; // CH=1 OP=3
cfg[1530] = { 1'b0, 8'h52, 8'h15}; // CH=2 OP=0
cfg[1531] = { 1'b1, 8'h83, 8'h73}; // CH=6 OP=0
cfg[1532] = { 1'b0, 8'h52, 8'ha1}; // CH=2 OP=0
cfg[1533] = { 1'b1, 8'hcd, 8'h55}; // CH=4 OP=3
cfg[1534] = { 1'b1, 8'h46, 8'h9e}; // CH=5 OP=1
cfg[1535] = { 1'b0, 8'h56, 8'hbd}; // CH=2 OP=1
cfg[1536] = { 1'b1, 8'h7a, 8'he8}; // CH=5 OP=2
cfg[1537] = { 1'b1, 8'hf1, 8'hac}; // CH=4 OP=0
cfg[1538] = { 1'b1, 8'hb9, 8'hd8}; // CH=4 OP=2
cfg[1539] = { 1'b0, 8'hbd, 8'h96}; // CH=1 OP=3
cfg[1540] = { 1'b1, 8'hd2, 8'h75}; // CH=5 OP=0
cfg[1541] = { 1'b0, 8'h45, 8'h76}; // CH=1 OP=1
cfg[1542] = { 1'b1, 8'he7, 8'h1a}; // CH=6 OP=1
cfg[1543] = { 1'b1, 8'h3c, 8'hab}; // CH=3 OP=3
cfg[1544] = { 1'b0, 8'hda, 8'hba}; // CH=2 OP=2
cfg[1545] = { 1'b1, 8'h97, 8'h93}; // CH=6 OP=1
cfg[1546] = { 1'b1, 8'h7f, 8'h20}; // CH=6 OP=3
cfg[1547] = { 1'b1, 8'h48, 8'h61}; // CH=3 OP=2
cfg[1548] = { 1'b0, 8'he9, 8'h4}; // CH=1 OP=2
cfg[1549] = { 1'b0, 8'h34, 8'hbf}; // CH=0 OP=1
cfg[1550] = { 1'b1, 8'hd2, 8'h91}; // CH=5 OP=0
cfg[1551] = { 1'b1, 8'hf4, 8'hd7}; // CH=3 OP=1
cfg[1552] = { 1'b1, 8'h67, 8'hbe}; // CH=6 OP=1
cfg[1553] = { 1'b1, 8'ha8, 8'hfa}; // CH=3 OP=2
cfg[1554] = { 1'b1, 8'h98, 8'hd4}; // CH=3 OP=2
cfg[1555] = { 1'b1, 8'hb9, 8'hc}; // CH=4 OP=2
cfg[1556] = { 1'b1, 8'hac, 8'h64}; // CH=3 OP=3
cfg[1557] = { 1'b1, 8'hae, 8'h1a}; // CH=5 OP=3
cfg[1558] = { 1'b0, 8'h6d, 8'hb5}; // CH=1 OP=3
cfg[1559] = { 1'b0, 8'hff, 8'hc4}; // CH=3 OP=3
cfg[1560] = { 1'b1, 8'hd6, 8'h4a}; // CH=5 OP=1
cfg[1561] = { 1'b1, 8'h94, 8'he9}; // CH=3 OP=1
cfg[1562] = { 1'b0, 8'h8e, 8'h34}; // CH=2 OP=3
cfg[1563] = { 1'b0, 8'h62, 8'h3a}; // CH=2 OP=0
cfg[1564] = { 1'b1, 8'hcd, 8'hd2}; // CH=4 OP=3
cfg[1565] = { 1'b0, 8'hb8, 8'h8b}; // CH=0 OP=2
cfg[1566] = { 1'b0, 8'hcf, 8'ha6}; // CH=3 OP=3
cfg[1567] = { 1'b0, 8'he9, 8'hbb}; // CH=1 OP=2
cfg[1568] = { 1'b1, 8'h9e, 8'hb9}; // CH=5 OP=3
cfg[1569] = { 1'b0, 8'h63, 8'heb}; // CH=3 OP=0
cfg[1570] = { 1'b1, 8'had, 8'hf0}; // CH=4 OP=3
cfg[1571] = { 1'b1, 8'h96, 8'he9}; // CH=5 OP=1
cfg[1572] = { 1'b1, 8'hcb, 8'h4a}; // CH=6 OP=2
cfg[1573] = { 1'b1, 8'hc9, 8'h52}; // CH=4 OP=2
cfg[1574] = { 1'b0, 8'h97, 8'hd7}; // CH=3 OP=1
cfg[1575] = { 1'b0, 8'h4f, 8'h63}; // CH=3 OP=3
cfg[1576] = { 1'b0, 8'hca, 8'h9}; // CH=2 OP=2
cfg[1577] = { 1'b0, 8'hcd, 8'h8}; // CH=1 OP=3
cfg[1578] = { 1'b1, 8'h3e, 8'ha6}; // CH=5 OP=3
cfg[1579] = { 1'b0, 8'had, 8'h9}; // CH=1 OP=3
cfg[1580] = { 1'b1, 8'hf3, 8'hb6}; // CH=6 OP=0
cfg[1581] = { 1'b0, 8'hcc, 8'h4d}; // CH=0 OP=3
cfg[1582] = { 1'b0, 8'h34, 8'h18}; // CH=0 OP=1
cfg[1583] = { 1'b1, 8'hfd, 8'h1d}; // CH=4 OP=3
cfg[1584] = { 1'b1, 8'h94, 8'hf4}; // CH=3 OP=1
cfg[1585] = { 1'b1, 8'he4, 8'h57}; // CH=3 OP=1
cfg[1586] = { 1'b1, 8'h77, 8'h60}; // CH=6 OP=1
cfg[1587] = { 1'b0, 8'h45, 8'ha}; // CH=1 OP=1
cfg[1588] = { 1'b1, 8'h83, 8'hb1}; // CH=6 OP=0
cfg[1589] = { 1'b0, 8'h30, 8'hba}; // CH=0 OP=0
cfg[1590] = { 1'b1, 8'ha5, 8'h71}; // CH=4 OP=1
cfg[1591] = { 1'b0, 8'h32, 8'hf0}; // CH=2 OP=0
cfg[1592] = { 1'b0, 8'hf3, 8'h24}; // CH=3 OP=0
cfg[1593] = { 1'b1, 8'he7, 8'h7a}; // CH=6 OP=1
cfg[1594] = { 1'b0, 8'h3f, 8'hb1}; // CH=3 OP=3
cfg[1595] = { 1'b0, 8'h9f, 8'h5e}; // CH=3 OP=3
cfg[1596] = { 1'b0, 8'hc4, 8'hd5}; // CH=0 OP=1
cfg[1597] = { 1'b1, 8'h65, 8'h1a}; // CH=4 OP=1
cfg[1598] = { 1'b0, 8'h6f, 8'h9d}; // CH=3 OP=3
cfg[1599] = { 1'b0, 8'hd2, 8'hce}; // CH=2 OP=0
cfg[1600] = { 1'b1, 8'h78, 8'hf1}; // CH=3 OP=2
cfg[1601] = { 1'b1, 8'haa, 8'he1}; // CH=5 OP=2
cfg[1602] = { 1'b1, 8'hbb, 8'h5}; // CH=6 OP=2
cfg[1603] = { 1'b0, 8'h35, 8'h27}; // CH=1 OP=1
cfg[1604] = { 1'b0, 8'he6, 8'hdd}; // CH=2 OP=1
cfg[1605] = { 1'b1, 8'h44, 8'h77}; // CH=3 OP=1
cfg[1606] = { 1'b0, 8'h94, 8'h13}; // CH=0 OP=1
cfg[1607] = { 1'b0, 8'hfa, 8'h34}; // CH=2 OP=2
cfg[1608] = { 1'b0, 8'h69, 8'hd1}; // CH=1 OP=2
cfg[1609] = { 1'b1, 8'h3c, 8'h9f}; // CH=3 OP=3
cfg[1610] = { 1'b0, 8'hb4, 8'h91}; // CH=0 OP=1
cfg[1611] = { 1'b0, 8'h5e, 8'h72}; // CH=2 OP=3
cfg[1612] = { 1'b1, 8'h9f, 8'h78}; // CH=6 OP=3
cfg[1613] = { 1'b0, 8'h7c, 8'hfe}; // CH=0 OP=3
cfg[1614] = { 1'b0, 8'hf3, 8'h2f}; // CH=3 OP=0
cfg[1615] = { 1'b0, 8'h91, 8'hff}; // CH=1 OP=0
cfg[1616] = { 1'b0, 8'hc5, 8'hc1}; // CH=1 OP=1
cfg[1617] = { 1'b0, 8'h97, 8'hd3}; // CH=3 OP=1
cfg[1618] = { 1'b1, 8'h36, 8'hf8}; // CH=5 OP=1
cfg[1619] = { 1'b1, 8'hc7, 8'ha1}; // CH=6 OP=1
cfg[1620] = { 1'b1, 8'h3a, 8'h8b}; // CH=5 OP=2
cfg[1621] = { 1'b1, 8'hb2, 8'h8c}; // CH=5 OP=0
cfg[1622] = { 1'b0, 8'h51, 8'h98}; // CH=1 OP=0
cfg[1623] = { 1'b0, 8'hcd, 8'h96}; // CH=1 OP=3
cfg[1624] = { 1'b0, 8'hc0, 8'hc5}; // CH=0 OP=0
cfg[1625] = { 1'b0, 8'hc6, 8'hc5}; // CH=2 OP=1
cfg[1626] = { 1'b0, 8'h87, 8'h59}; // CH=3 OP=1
cfg[1627] = { 1'b1, 8'h5b, 8'he7}; // CH=6 OP=2
cfg[1628] = { 1'b0, 8'h53, 8'hde}; // CH=3 OP=0
cfg[1629] = { 1'b1, 8'hf4, 8'h12}; // CH=3 OP=1
cfg[1630] = { 1'b0, 8'h7f, 8'hf9}; // CH=3 OP=3
cfg[1631] = { 1'b0, 8'h30, 8'h3f}; // CH=0 OP=0
cfg[1632] = { 1'b1, 8'h81, 8'ha4}; // CH=4 OP=0
cfg[1633] = { 1'b0, 8'h4e, 8'h3b}; // CH=2 OP=3
cfg[1634] = { 1'b0, 8'h83, 8'h0}; // CH=3 OP=0
cfg[1635] = { 1'b1, 8'h6d, 8'hd5}; // CH=4 OP=3
cfg[1636] = { 1'b0, 8'hb7, 8'h5c}; // CH=3 OP=1
cfg[1637] = { 1'b1, 8'he0, 8'he4}; // CH=3 OP=0
cfg[1638] = { 1'b0, 8'hef, 8'hff}; // CH=3 OP=3
cfg[1639] = { 1'b1, 8'h8b, 8'ha3}; // CH=6 OP=2
cfg[1640] = { 1'b1, 8'h55, 8'hcc}; // CH=4 OP=1
cfg[1641] = { 1'b0, 8'ha3, 8'h6a}; // CH=3 OP=0
cfg[1642] = { 1'b0, 8'hb2, 8'h6b}; // CH=2 OP=0
cfg[1643] = { 1'b1, 8'h87, 8'h30}; // CH=6 OP=1
cfg[1644] = { 1'b0, 8'he3, 8'h4f}; // CH=3 OP=0
cfg[1645] = { 1'b1, 8'h9b, 8'h54}; // CH=6 OP=2
cfg[1646] = { 1'b0, 8'ha6, 8'h38}; // CH=2 OP=1
cfg[1647] = { 1'b0, 8'ha5, 8'h2e}; // CH=1 OP=1
cfg[1648] = { 1'b0, 8'h57, 8'h1e}; // CH=3 OP=1
cfg[1649] = { 1'b0, 8'hdf, 8'haf}; // CH=3 OP=3
cfg[1650] = { 1'b0, 8'h49, 8'h2e}; // CH=1 OP=2
cfg[1651] = { 1'b1, 8'hb4, 8'h6f}; // CH=3 OP=1
cfg[1652] = { 1'b1, 8'he5, 8'h32}; // CH=4 OP=1
cfg[1653] = { 1'b0, 8'h34, 8'h63}; // CH=0 OP=1
cfg[1654] = { 1'b0, 8'h88, 8'hb0}; // CH=0 OP=2
cfg[1655] = { 1'b1, 8'hc1, 8'h60}; // CH=4 OP=0
cfg[1656] = { 1'b1, 8'hef, 8'hf0}; // CH=6 OP=3
cfg[1657] = { 1'b0, 8'h4b, 8'ha4}; // CH=3 OP=2
cfg[1658] = { 1'b0, 8'hfa, 8'h5a}; // CH=2 OP=2
cfg[1659] = { 1'b1, 8'hd9, 8'h72}; // CH=4 OP=2
cfg[1660] = { 1'b1, 8'hca, 8'ha1}; // CH=5 OP=2
cfg[1661] = { 1'b0, 8'ha0, 8'hd7}; // CH=0 OP=0
cfg[1662] = { 1'b0, 8'hfc, 8'hbc}; // CH=0 OP=3
cfg[1663] = { 1'b1, 8'h3c, 8'hf0}; // CH=3 OP=3
cfg[1664] = { 1'b1, 8'hb5, 8'h79}; // CH=4 OP=1
cfg[1665] = { 1'b0, 8'ha5, 8'h98}; // CH=1 OP=1
cfg[1666] = { 1'b1, 8'h4a, 8'hbf}; // CH=5 OP=2
cfg[1667] = { 1'b1, 8'h46, 8'ha}; // CH=5 OP=1
cfg[1668] = { 1'b1, 8'h6d, 8'h4}; // CH=4 OP=3
cfg[1669] = { 1'b1, 8'ha4, 8'hde}; // CH=3 OP=1
cfg[1670] = { 1'b1, 8'hb4, 8'hde}; // CH=3 OP=1
cfg[1671] = { 1'b0, 8'hf7, 8'h7e}; // CH=3 OP=1
cfg[1672] = { 1'b1, 8'h9c, 8'h7b}; // CH=3 OP=3
cfg[1673] = { 1'b1, 8'hf2, 8'hb7}; // CH=5 OP=0
cfg[1674] = { 1'b0, 8'ha7, 8'hcf}; // CH=3 OP=1
cfg[1675] = { 1'b0, 8'h4d, 8'h67}; // CH=1 OP=3
cfg[1676] = { 1'b0, 8'h97, 8'h26}; // CH=3 OP=1
cfg[1677] = { 1'b1, 8'hdd, 8'h30}; // CH=4 OP=3
cfg[1678] = { 1'b0, 8'h4a, 8'h35}; // CH=2 OP=2
cfg[1679] = { 1'b1, 8'h5e, 8'h13}; // CH=5 OP=3
cfg[1680] = { 1'b0, 8'h3c, 8'h14}; // CH=0 OP=3
cfg[1681] = { 1'b0, 8'hbb, 8'hec}; // CH=3 OP=2
cfg[1682] = { 1'b1, 8'h36, 8'h81}; // CH=5 OP=1
cfg[1683] = { 1'b0, 8'hed, 8'h7}; // CH=1 OP=3
cfg[1684] = { 1'b0, 8'hbc, 8'h5}; // CH=0 OP=3
cfg[1685] = { 1'b1, 8'ha0, 8'h3e}; // CH=3 OP=0
cfg[1686] = { 1'b0, 8'h39, 8'h97}; // CH=1 OP=2
cfg[1687] = { 1'b1, 8'h63, 8'h74}; // CH=6 OP=0
cfg[1688] = { 1'b0, 8'h90, 8'hbe}; // CH=0 OP=0
cfg[1689] = { 1'b1, 8'h62, 8'h1c}; // CH=5 OP=0
cfg[1690] = { 1'b1, 8'he9, 8'h59}; // CH=4 OP=2
cfg[1691] = { 1'b1, 8'h66, 8'h14}; // CH=5 OP=1
cfg[1692] = { 1'b1, 8'h80, 8'h4a}; // CH=3 OP=0
cfg[1693] = { 1'b0, 8'h8c, 8'h37}; // CH=0 OP=3
cfg[1694] = { 1'b1, 8'h40, 8'hf4}; // CH=3 OP=0
cfg[1695] = { 1'b1, 8'h40, 8'h18}; // CH=3 OP=0
cfg[1696] = { 1'b1, 8'hd8, 8'h62}; // CH=3 OP=2
cfg[1697] = { 1'b0, 8'h4c, 8'hdd}; // CH=0 OP=3
cfg[1698] = { 1'b1, 8'h5c, 8'h8d}; // CH=3 OP=3
cfg[1699] = { 1'b0, 8'hbe, 8'h27}; // CH=2 OP=3
cfg[1700] = { 1'b1, 8'ha7, 8'h80}; // CH=6 OP=1
cfg[1701] = { 1'b1, 8'h30, 8'h94}; // CH=3 OP=0
cfg[1702] = { 1'b0, 8'h7c, 8'h8e}; // CH=0 OP=3
cfg[1703] = { 1'b0, 8'hcd, 8'h1b}; // CH=1 OP=3
cfg[1704] = { 1'b0, 8'h5d, 8'h5b}; // CH=1 OP=3
cfg[1705] = { 1'b0, 8'h8c, 8'h9b}; // CH=0 OP=3
cfg[1706] = { 1'b0, 8'hf5, 8'h73}; // CH=1 OP=1
cfg[1707] = { 1'b0, 8'hc0, 8'hc0}; // CH=0 OP=0
cfg[1708] = { 1'b1, 8'h40, 8'hcb}; // CH=3 OP=0
cfg[1709] = { 1'b0, 8'h67, 8'hdb}; // CH=3 OP=1
cfg[1710] = { 1'b1, 8'h52, 8'h82}; // CH=5 OP=0
cfg[1711] = { 1'b1, 8'h82, 8'h90}; // CH=5 OP=0
cfg[1712] = { 1'b0, 8'hfe, 8'h1f}; // CH=2 OP=3
cfg[1713] = { 1'b0, 8'hcc, 8'h3a}; // CH=0 OP=3
cfg[1714] = { 1'b0, 8'h30, 8'h95}; // CH=0 OP=0
cfg[1715] = { 1'b1, 8'ha4, 8'hac}; // CH=3 OP=1
cfg[1716] = { 1'b0, 8'h64, 8'he}; // CH=0 OP=1
cfg[1717] = { 1'b1, 8'h87, 8'hfe}; // CH=6 OP=1
cfg[1718] = { 1'b0, 8'h62, 8'h21}; // CH=2 OP=0
cfg[1719] = { 1'b1, 8'he5, 8'h94}; // CH=4 OP=1
cfg[1720] = { 1'b0, 8'h75, 8'h9c}; // CH=1 OP=1
cfg[1721] = { 1'b0, 8'h94, 8'h82}; // CH=0 OP=1
cfg[1722] = { 1'b1, 8'hce, 8'h7e}; // CH=5 OP=3
cfg[1723] = { 1'b1, 8'h63, 8'h84}; // CH=6 OP=0
cfg[1724] = { 1'b0, 8'h94, 8'hac}; // CH=0 OP=1
cfg[1725] = { 1'b1, 8'h38, 8'h58}; // CH=3 OP=2
cfg[1726] = { 1'b0, 8'h9c, 8'h67}; // CH=0 OP=3
cfg[1727] = { 1'b1, 8'hcb, 8'h65}; // CH=6 OP=2
cfg[1728] = { 1'b0, 8'hec, 8'ha3}; // CH=0 OP=3
cfg[1729] = { 1'b1, 8'h81, 8'h48}; // CH=4 OP=0
cfg[1730] = { 1'b0, 8'h7d, 8'h40}; // CH=1 OP=3
cfg[1731] = { 1'b1, 8'h34, 8'h9f}; // CH=3 OP=1
cfg[1732] = { 1'b1, 8'h79, 8'he0}; // CH=4 OP=2
cfg[1733] = { 1'b1, 8'he7, 8'h44}; // CH=6 OP=1
cfg[1734] = { 1'b1, 8'ha5, 8'hd8}; // CH=4 OP=1
cfg[1735] = { 1'b0, 8'hac, 8'hd8}; // CH=0 OP=3
cfg[1736] = { 1'b1, 8'h77, 8'h71}; // CH=6 OP=1
cfg[1737] = { 1'b0, 8'h63, 8'h14}; // CH=3 OP=0
cfg[1738] = { 1'b1, 8'he4, 8'h5d}; // CH=3 OP=1
cfg[1739] = { 1'b1, 8'h7a, 8'h9d}; // CH=5 OP=2
cfg[1740] = { 1'b0, 8'h8c, 8'ha0}; // CH=0 OP=3
cfg[1741] = { 1'b0, 8'h6d, 8'hbd}; // CH=1 OP=3
cfg[1742] = { 1'b1, 8'hb1, 8'h5e}; // CH=4 OP=0
cfg[1743] = { 1'b0, 8'h89, 8'hab}; // CH=1 OP=2
cfg[1744] = { 1'b1, 8'h99, 8'h51}; // CH=4 OP=2
cfg[1745] = { 1'b1, 8'h45, 8'h5d}; // CH=4 OP=1
cfg[1746] = { 1'b1, 8'hbc, 8'hcf}; // CH=3 OP=3
cfg[1747] = { 1'b1, 8'ha8, 8'he3}; // CH=3 OP=2
cfg[1748] = { 1'b0, 8'ha5, 8'h4}; // CH=1 OP=1
cfg[1749] = { 1'b0, 8'h36, 8'h5}; // CH=2 OP=1
cfg[1750] = { 1'b0, 8'hc3, 8'hac}; // CH=3 OP=0
cfg[1751] = { 1'b1, 8'hc8, 8'h19}; // CH=3 OP=2
cfg[1752] = { 1'b0, 8'hb5, 8'hca}; // CH=1 OP=1
cfg[1753] = { 1'b1, 8'hac, 8'h53}; // CH=3 OP=3
cfg[1754] = { 1'b0, 8'h7b, 8'hec}; // CH=3 OP=2
cfg[1755] = { 1'b0, 8'h5c, 8'h31}; // CH=0 OP=3
cfg[1756] = { 1'b1, 8'hce, 8'hed}; // CH=5 OP=3
cfg[1757] = { 1'b0, 8'h5c, 8'hb7}; // CH=0 OP=3
cfg[1758] = { 1'b1, 8'h7c, 8'h16}; // CH=3 OP=3
cfg[1759] = { 1'b1, 8'he6, 8'hbc}; // CH=5 OP=1
cfg[1760] = { 1'b1, 8'haf, 8'h41}; // CH=6 OP=3
cfg[1761] = { 1'b1, 8'h64, 8'hb}; // CH=3 OP=1
cfg[1762] = { 1'b1, 8'h4a, 8'h5e}; // CH=5 OP=2
cfg[1763] = { 1'b1, 8'h7b, 8'h29}; // CH=6 OP=2
cfg[1764] = { 1'b0, 8'h68, 8'h14}; // CH=0 OP=2
cfg[1765] = { 1'b1, 8'h74, 8'he3}; // CH=3 OP=1
cfg[1766] = { 1'b1, 8'h85, 8'hf2}; // CH=4 OP=1
cfg[1767] = { 1'b1, 8'h9b, 8'hdf}; // CH=6 OP=2
cfg[1768] = { 1'b1, 8'h57, 8'h2}; // CH=6 OP=1
cfg[1769] = { 1'b1, 8'h76, 8'he9}; // CH=5 OP=1
cfg[1770] = { 1'b0, 8'h58, 8'h98}; // CH=0 OP=2
cfg[1771] = { 1'b1, 8'ha7, 8'hfc}; // CH=6 OP=1
cfg[1772] = { 1'b1, 8'hb4, 8'hc}; // CH=3 OP=1
cfg[1773] = { 1'b1, 8'hde, 8'h97}; // CH=5 OP=3
cfg[1774] = { 1'b0, 8'hf2, 8'h7f}; // CH=2 OP=0
cfg[1775] = { 1'b0, 8'hd5, 8'h77}; // CH=1 OP=1
cfg[1776] = { 1'b1, 8'hc7, 8'h26}; // CH=6 OP=1
cfg[1777] = { 1'b0, 8'ha6, 8'h31}; // CH=2 OP=1
cfg[1778] = { 1'b1, 8'ha9, 8'hb9}; // CH=4 OP=2
cfg[1779] = { 1'b0, 8'h92, 8'h68}; // CH=2 OP=0
cfg[1780] = { 1'b0, 8'h40, 8'h59}; // CH=0 OP=0
cfg[1781] = { 1'b0, 8'he7, 8'h26}; // CH=3 OP=1
cfg[1782] = { 1'b0, 8'h9c, 8'h32}; // CH=0 OP=3
cfg[1783] = { 1'b1, 8'h7a, 8'hc9}; // CH=5 OP=2
cfg[1784] = { 1'b0, 8'h6c, 8'h49}; // CH=0 OP=3
cfg[1785] = { 1'b0, 8'h42, 8'hc0}; // CH=2 OP=0
cfg[1786] = { 1'b1, 8'h71, 8'he6}; // CH=4 OP=0
cfg[1787] = { 1'b1, 8'h8c, 8'hb0}; // CH=3 OP=3
cfg[1788] = { 1'b0, 8'hfe, 8'h59}; // CH=2 OP=3
cfg[1789] = { 1'b1, 8'he7, 8'heb}; // CH=6 OP=1
cfg[1790] = { 1'b0, 8'he6, 8'h15}; // CH=2 OP=1
cfg[1791] = { 1'b1, 8'h94, 8'hf}; // CH=3 OP=1
cfg[1792] = { 1'b1, 8'he6, 8'hab}; // CH=5 OP=1
cfg[1793] = { 1'b0, 8'h56, 8'h25}; // CH=2 OP=1
cfg[1794] = { 1'b1, 8'h4c, 8'h91}; // CH=3 OP=3
cfg[1795] = { 1'b1, 8'h3e, 8'hd3}; // CH=5 OP=3
cfg[1796] = { 1'b1, 8'haf, 8'hdd}; // CH=6 OP=3
cfg[1797] = { 1'b1, 8'h3c, 8'h8d}; // CH=3 OP=3
cfg[1798] = { 1'b1, 8'h3a, 8'he6}; // CH=5 OP=2
cfg[1799] = { 1'b0, 8'hd8, 8'hd1}; // CH=0 OP=2
cfg[1800] = { 1'b0, 8'hbf, 8'h49}; // CH=3 OP=3
cfg[1801] = { 1'b1, 8'h53, 8'h58}; // CH=6 OP=0
cfg[1802] = { 1'b0, 8'h39, 8'h3}; // CH=1 OP=2
cfg[1803] = { 1'b0, 8'h8f, 8'h28}; // CH=3 OP=3
cfg[1804] = { 1'b0, 8'hdc, 8'hb9}; // CH=0 OP=3
cfg[1805] = { 1'b1, 8'ha9, 8'h8d}; // CH=4 OP=2
cfg[1806] = { 1'b0, 8'he6, 8'hc9}; // CH=2 OP=1
cfg[1807] = { 1'b1, 8'hf3, 8'h5}; // CH=6 OP=0
cfg[1808] = { 1'b1, 8'h3a, 8'h40}; // CH=5 OP=2
cfg[1809] = { 1'b0, 8'h94, 8'h61}; // CH=0 OP=1
cfg[1810] = { 1'b0, 8'hb5, 8'hd1}; // CH=1 OP=1
cfg[1811] = { 1'b0, 8'h43, 8'h25}; // CH=3 OP=0
cfg[1812] = { 1'b1, 8'hee, 8'h5e}; // CH=5 OP=3
cfg[1813] = { 1'b1, 8'hca, 8'he7}; // CH=5 OP=2
cfg[1814] = { 1'b1, 8'he4, 8'h74}; // CH=3 OP=1
cfg[1815] = { 1'b0, 8'had, 8'hde}; // CH=1 OP=3
cfg[1816] = { 1'b0, 8'hb3, 8'hd5}; // CH=3 OP=0
cfg[1817] = { 1'b1, 8'hf3, 8'hb2}; // CH=6 OP=0
cfg[1818] = { 1'b1, 8'h54, 8'h60}; // CH=3 OP=1
cfg[1819] = { 1'b0, 8'hff, 8'hf4}; // CH=3 OP=3
cfg[1820] = { 1'b1, 8'h94, 8'ha9}; // CH=3 OP=1
cfg[1821] = { 1'b0, 8'hf3, 8'h7}; // CH=3 OP=0
cfg[1822] = { 1'b1, 8'he1, 8'h34}; // CH=4 OP=0
cfg[1823] = { 1'b1, 8'hab, 8'h1b}; // CH=6 OP=2
cfg[1824] = { 1'b0, 8'h8f, 8'h8f}; // CH=3 OP=3
cfg[1825] = { 1'b0, 8'h3c, 8'h6d}; // CH=0 OP=3
cfg[1826] = { 1'b0, 8'hef, 8'h42}; // CH=3 OP=3
cfg[1827] = { 1'b1, 8'he2, 8'hf4}; // CH=5 OP=0
cfg[1828] = { 1'b1, 8'h37, 8'h54}; // CH=6 OP=1
cfg[1829] = { 1'b1, 8'h36, 8'h48}; // CH=5 OP=1
cfg[1830] = { 1'b0, 8'h37, 8'hf1}; // CH=3 OP=1
cfg[1831] = { 1'b1, 8'h3e, 8'hdd}; // CH=5 OP=3
cfg[1832] = { 1'b0, 8'h73, 8'hd1}; // CH=3 OP=0
cfg[1833] = { 1'b1, 8'h8e, 8'h10}; // CH=5 OP=3
cfg[1834] = { 1'b0, 8'h71, 8'h1e}; // CH=1 OP=0
cfg[1835] = { 1'b0, 8'had, 8'h8b}; // CH=1 OP=3
cfg[1836] = { 1'b0, 8'h9d, 8'hce}; // CH=1 OP=3
cfg[1837] = { 1'b1, 8'h7f, 8'hc2}; // CH=6 OP=3
cfg[1838] = { 1'b0, 8'hb6, 8'h17}; // CH=2 OP=1
cfg[1839] = { 1'b1, 8'hec, 8'h5f}; // CH=3 OP=3
cfg[1840] = { 1'b0, 8'h62, 8'h51}; // CH=2 OP=0
cfg[1841] = { 1'b1, 8'hd5, 8'hff}; // CH=4 OP=1
cfg[1842] = { 1'b0, 8'h64, 8'hf}; // CH=0 OP=1
cfg[1843] = { 1'b0, 8'h82, 8'h2d}; // CH=2 OP=0
cfg[1844] = { 1'b1, 8'h9c, 8'hd1}; // CH=3 OP=3
cfg[1845] = { 1'b1, 8'h39, 8'hdb}; // CH=4 OP=2
cfg[1846] = { 1'b1, 8'hb9, 8'h9e}; // CH=4 OP=2
cfg[1847] = { 1'b1, 8'h6f, 8'hb5}; // CH=6 OP=3
cfg[1848] = { 1'b1, 8'h5c, 8'h14}; // CH=3 OP=3
cfg[1849] = { 1'b1, 8'h80, 8'h65}; // CH=3 OP=0
cfg[1850] = { 1'b0, 8'he2, 8'h94}; // CH=2 OP=0
cfg[1851] = { 1'b1, 8'hb8, 8'h93}; // CH=3 OP=2
cfg[1852] = { 1'b1, 8'had, 8'ha3}; // CH=4 OP=3
cfg[1853] = { 1'b0, 8'h9c, 8'h9e}; // CH=0 OP=3
cfg[1854] = { 1'b0, 8'h38, 8'hab}; // CH=0 OP=2
cfg[1855] = { 1'b1, 8'h72, 8'h87}; // CH=5 OP=0
cfg[1856] = { 1'b0, 8'ha8, 8'h25}; // CH=0 OP=2
cfg[1857] = { 1'b0, 8'hee, 8'h9a}; // CH=2 OP=3
cfg[1858] = { 1'b0, 8'h54, 8'h3a}; // CH=0 OP=1
cfg[1859] = { 1'b0, 8'he8, 8'h68}; // CH=0 OP=2
cfg[1860] = { 1'b1, 8'h7b, 8'hfb}; // CH=6 OP=2
cfg[1861] = { 1'b1, 8'hd7, 8'h2a}; // CH=6 OP=1
cfg[1862] = { 1'b1, 8'h73, 8'hcb}; // CH=6 OP=0
cfg[1863] = { 1'b1, 8'hab, 8'h76}; // CH=6 OP=2
cfg[1864] = { 1'b0, 8'h9f, 8'hfd}; // CH=3 OP=3
cfg[1865] = { 1'b0, 8'h47, 8'h48}; // CH=3 OP=1
cfg[1866] = { 1'b0, 8'h62, 8'he3}; // CH=2 OP=0
cfg[1867] = { 1'b1, 8'h9c, 8'hd9}; // CH=3 OP=3
cfg[1868] = { 1'b1, 8'ha9, 8'h50}; // CH=4 OP=2
cfg[1869] = { 1'b1, 8'hba, 8'ha2}; // CH=5 OP=2
cfg[1870] = { 1'b1, 8'he7, 8'hc1}; // CH=6 OP=1
cfg[1871] = { 1'b0, 8'hb2, 8'hb0}; // CH=2 OP=0
cfg[1872] = { 1'b1, 8'hcd, 8'h41}; // CH=4 OP=3
cfg[1873] = { 1'b0, 8'h6c, 8'h3c}; // CH=0 OP=3
cfg[1874] = { 1'b0, 8'hb3, 8'h84}; // CH=3 OP=0
cfg[1875] = { 1'b1, 8'h30, 8'h67}; // CH=3 OP=0
cfg[1876] = { 1'b1, 8'h6f, 8'hb1}; // CH=6 OP=3
cfg[1877] = { 1'b1, 8'h96, 8'hb5}; // CH=5 OP=1
cfg[1878] = { 1'b0, 8'h38, 8'hb4}; // CH=0 OP=2
cfg[1879] = { 1'b0, 8'hf9, 8'hdd}; // CH=1 OP=2
cfg[1880] = { 1'b1, 8'ha9, 8'hdd}; // CH=4 OP=2
cfg[1881] = { 1'b1, 8'hea, 8'h50}; // CH=5 OP=2
cfg[1882] = { 1'b1, 8'hb8, 8'h6f}; // CH=3 OP=2
cfg[1883] = { 1'b1, 8'hd8, 8'hab}; // CH=3 OP=2
cfg[1884] = { 1'b1, 8'hed, 8'h97}; // CH=4 OP=3
cfg[1885] = { 1'b1, 8'h9f, 8'hd8}; // CH=6 OP=3
cfg[1886] = { 1'b0, 8'h54, 8'h69}; // CH=0 OP=1
cfg[1887] = { 1'b0, 8'hd6, 8'ha3}; // CH=2 OP=1
cfg[1888] = { 1'b1, 8'hd0, 8'he6}; // CH=3 OP=0
cfg[1889] = { 1'b0, 8'h79, 8'hc4}; // CH=1 OP=2
cfg[1890] = { 1'b1, 8'h64, 8'h14}; // CH=3 OP=1
cfg[1891] = { 1'b0, 8'h90, 8'h83}; // CH=0 OP=0
cfg[1892] = { 1'b0, 8'hb4, 8'h40}; // CH=0 OP=1
cfg[1893] = { 1'b0, 8'hf5, 8'h18}; // CH=1 OP=1
cfg[1894] = { 1'b0, 8'hcd, 8'hb6}; // CH=1 OP=3
cfg[1895] = { 1'b1, 8'h36, 8'hbe}; // CH=5 OP=1
cfg[1896] = { 1'b1, 8'hd9, 8'h5c}; // CH=4 OP=2
cfg[1897] = { 1'b0, 8'h70, 8'h32}; // CH=0 OP=0
cfg[1898] = { 1'b1, 8'he2, 8'h2}; // CH=5 OP=0
cfg[1899] = { 1'b1, 8'he1, 8'h7c}; // CH=4 OP=0
cfg[1900] = { 1'b1, 8'h95, 8'he0}; // CH=4 OP=1
cfg[1901] = { 1'b1, 8'h73, 8'hfc}; // CH=6 OP=0
cfg[1902] = { 1'b0, 8'hd1, 8'hd9}; // CH=1 OP=0
cfg[1903] = { 1'b1, 8'hc6, 8'hf6}; // CH=5 OP=1
cfg[1904] = { 1'b1, 8'h93, 8'hac}; // CH=6 OP=0
cfg[1905] = { 1'b0, 8'hc9, 8'h6a}; // CH=1 OP=2
cfg[1906] = { 1'b1, 8'ha2, 8'hc6}; // CH=5 OP=0
cfg[1907] = { 1'b0, 8'he5, 8'hf9}; // CH=1 OP=1
cfg[1908] = { 1'b1, 8'h92, 8'hf4}; // CH=5 OP=0
cfg[1909] = { 1'b1, 8'h53, 8'hd5}; // CH=6 OP=0
cfg[1910] = { 1'b1, 8'h98, 8'h6b}; // CH=3 OP=2
cfg[1911] = { 1'b1, 8'h90, 8'h90}; // CH=3 OP=0
cfg[1912] = { 1'b0, 8'he5, 8'hdd}; // CH=1 OP=1
cfg[1913] = { 1'b0, 8'h40, 8'ha4}; // CH=0 OP=0
cfg[1914] = { 1'b1, 8'h40, 8'h37}; // CH=3 OP=0
cfg[1915] = { 1'b1, 8'h39, 8'h1}; // CH=4 OP=2
cfg[1916] = { 1'b0, 8'h35, 8'ha3}; // CH=1 OP=1
cfg[1917] = { 1'b1, 8'h32, 8'hb6}; // CH=5 OP=0
cfg[1918] = { 1'b0, 8'haa, 8'hac}; // CH=2 OP=2
cfg[1919] = { 1'b0, 8'heb, 8'h0}; // CH=3 OP=2
cfg[1920] = { 1'b0, 8'h7b, 8'h55}; // CH=3 OP=2
cfg[1921] = { 1'b0, 8'he5, 8'he5}; // CH=1 OP=1
cfg[1922] = { 1'b0, 8'h46, 8'hca}; // CH=2 OP=1
cfg[1923] = { 1'b0, 8'h53, 8'ha}; // CH=3 OP=0
cfg[1924] = { 1'b1, 8'hca, 8'h4a}; // CH=5 OP=2
cfg[1925] = { 1'b0, 8'hb9, 8'h83}; // CH=1 OP=2
cfg[1926] = { 1'b1, 8'hd3, 8'hb8}; // CH=6 OP=0
cfg[1927] = { 1'b0, 8'h80, 8'h62}; // CH=0 OP=0
cfg[1928] = { 1'b0, 8'h80, 8'he2}; // CH=0 OP=0
cfg[1929] = { 1'b1, 8'h72, 8'hcd}; // CH=5 OP=0
cfg[1930] = { 1'b1, 8'h57, 8'hbd}; // CH=6 OP=1
cfg[1931] = { 1'b0, 8'h74, 8'h3f}; // CH=0 OP=1
cfg[1932] = { 1'b1, 8'hc7, 8'h2b}; // CH=6 OP=1
cfg[1933] = { 1'b0, 8'h92, 8'h75}; // CH=2 OP=0
cfg[1934] = { 1'b1, 8'h9a, 8'hf9}; // CH=5 OP=2
cfg[1935] = { 1'b1, 8'hda, 8'hb2}; // CH=5 OP=2
cfg[1936] = { 1'b1, 8'h4c, 8'h85}; // CH=3 OP=3
cfg[1937] = { 1'b1, 8'h68, 8'h5}; // CH=3 OP=2
cfg[1938] = { 1'b0, 8'h85, 8'h85}; // CH=1 OP=1
cfg[1939] = { 1'b1, 8'hf8, 8'h9e}; // CH=3 OP=2
cfg[1940] = { 1'b0, 8'h4f, 8'h5b}; // CH=3 OP=3
cfg[1941] = { 1'b1, 8'h71, 8'h9a}; // CH=4 OP=0
cfg[1942] = { 1'b1, 8'h9c, 8'hff}; // CH=3 OP=3
cfg[1943] = { 1'b1, 8'h33, 8'hc1}; // CH=6 OP=0
cfg[1944] = { 1'b0, 8'hcd, 8'hb}; // CH=1 OP=3
cfg[1945] = { 1'b1, 8'ha7, 8'hbd}; // CH=6 OP=1
cfg[1946] = { 1'b0, 8'hf3, 8'h42}; // CH=3 OP=0
cfg[1947] = { 1'b0, 8'h5b, 8'h48}; // CH=3 OP=2
cfg[1948] = { 1'b0, 8'he1, 8'hcd}; // CH=1 OP=0
cfg[1949] = { 1'b1, 8'hd9, 8'h6b}; // CH=4 OP=2
cfg[1950] = { 1'b0, 8'hc7, 8'hc6}; // CH=3 OP=1
cfg[1951] = { 1'b0, 8'ha0, 8'h99}; // CH=0 OP=0
cfg[1952] = { 1'b1, 8'h41, 8'h36}; // CH=4 OP=0
cfg[1953] = { 1'b1, 8'h74, 8'h48}; // CH=3 OP=1
cfg[1954] = { 1'b1, 8'h42, 8'h53}; // CH=5 OP=0
cfg[1955] = { 1'b1, 8'he9, 8'h10}; // CH=4 OP=2
cfg[1956] = { 1'b1, 8'hdd, 8'h52}; // CH=4 OP=3
cfg[1957] = { 1'b1, 8'h38, 8'h9a}; // CH=3 OP=2
cfg[1958] = { 1'b1, 8'h71, 8'h68}; // CH=4 OP=0
cfg[1959] = { 1'b1, 8'hd3, 8'hf2}; // CH=6 OP=0
cfg[1960] = { 1'b0, 8'h9a, 8'h1b}; // CH=2 OP=2
cfg[1961] = { 1'b0, 8'h3a, 8'hb4}; // CH=2 OP=2
cfg[1962] = { 1'b0, 8'h7c, 8'hea}; // CH=0 OP=3
cfg[1963] = { 1'b1, 8'hf0, 8'h32}; // CH=3 OP=0
cfg[1964] = { 1'b0, 8'h32, 8'h85}; // CH=2 OP=0
cfg[1965] = { 1'b1, 8'h71, 8'h95}; // CH=4 OP=0
cfg[1966] = { 1'b0, 8'h78, 8'hf9}; // CH=0 OP=2
cfg[1967] = { 1'b0, 8'hbe, 8'h31}; // CH=2 OP=3
cfg[1968] = { 1'b0, 8'hbe, 8'h4b}; // CH=2 OP=3
cfg[1969] = { 1'b1, 8'h58, 8'h2}; // CH=3 OP=2
cfg[1970] = { 1'b0, 8'h52, 8'h9c}; // CH=2 OP=0
cfg[1971] = { 1'b1, 8'hac, 8'hd6}; // CH=3 OP=3
cfg[1972] = { 1'b1, 8'h43, 8'h52}; // CH=6 OP=0
cfg[1973] = { 1'b0, 8'h75, 8'haf}; // CH=1 OP=1
cfg[1974] = { 1'b1, 8'h91, 8'h45}; // CH=4 OP=0
cfg[1975] = { 1'b0, 8'h8a, 8'h2d}; // CH=2 OP=2
cfg[1976] = { 1'b1, 8'hbc, 8'haf}; // CH=3 OP=3
cfg[1977] = { 1'b1, 8'h58, 8'h9a}; // CH=3 OP=2
cfg[1978] = { 1'b0, 8'hb0, 8'h6}; // CH=0 OP=0
cfg[1979] = { 1'b1, 8'haa, 8'ha2}; // CH=5 OP=2
cfg[1980] = { 1'b0, 8'ha1, 8'haf}; // CH=1 OP=0
cfg[1981] = { 1'b1, 8'hcb, 8'hd6}; // CH=6 OP=2
cfg[1982] = { 1'b0, 8'h7b, 8'h7c}; // CH=3 OP=2
cfg[1983] = { 1'b1, 8'hc0, 8'haa}; // CH=3 OP=0
cfg[1984] = { 1'b1, 8'hed, 8'h48}; // CH=4 OP=3
cfg[1985] = { 1'b1, 8'h9c, 8'h5f}; // CH=3 OP=3
cfg[1986] = { 1'b1, 8'h36, 8'h34}; // CH=5 OP=1
cfg[1987] = { 1'b0, 8'h8e, 8'h38}; // CH=2 OP=3
cfg[1988] = { 1'b1, 8'h3e, 8'h3e}; // CH=5 OP=3
cfg[1989] = { 1'b0, 8'h41, 8'he0}; // CH=1 OP=0
cfg[1990] = { 1'b0, 8'hf0, 8'h59}; // CH=0 OP=0
cfg[1991] = { 1'b1, 8'hc6, 8'h24}; // CH=5 OP=1
cfg[1992] = { 1'b1, 8'h43, 8'h32}; // CH=6 OP=0
cfg[1993] = { 1'b0, 8'hed, 8'hb5}; // CH=1 OP=3
cfg[1994] = { 1'b0, 8'h35, 8'hca}; // CH=1 OP=1
cfg[1995] = { 1'b1, 8'h95, 8'h6a}; // CH=4 OP=1
cfg[1996] = { 1'b1, 8'hc9, 8'hc5}; // CH=4 OP=2
cfg[1997] = { 1'b0, 8'he4, 8'h28}; // CH=0 OP=1
cfg[1998] = { 1'b1, 8'h64, 8'h40}; // CH=3 OP=1
cfg[1999] = { 1'b1, 8'h54, 8'h7a}; // CH=3 OP=1
cfg[2000] = { 1'b0, 8'heb, 8'h9e}; // CH=3 OP=2
cfg[2001] = { 1'b0, 8'hc1, 8'h5d}; // CH=1 OP=0
cfg[2002] = { 1'b1, 8'h57, 8'h4a}; // CH=6 OP=1
cfg[2003] = { 1'b0, 8'hda, 8'h80}; // CH=2 OP=2
cfg[2004] = { 1'b0, 8'hfa, 8'h15}; // CH=2 OP=2
cfg[2005] = { 1'b1, 8'h50, 8'hde}; // CH=3 OP=0
cfg[2006] = { 1'b1, 8'h34, 8'he0}; // CH=3 OP=1
cfg[2007] = { 1'b0, 8'h57, 8'h21}; // CH=3 OP=1
cfg[2008] = { 1'b1, 8'hbb, 8'h42}; // CH=6 OP=2
cfg[2009] = { 1'b0, 8'h5a, 8'hbc}; // CH=2 OP=2
cfg[2010] = { 1'b0, 8'h87, 8'h6}; // CH=3 OP=1
cfg[2011] = { 1'b0, 8'hd2, 8'haf}; // CH=2 OP=0
cfg[2012] = { 1'b1, 8'h52, 8'hff}; // CH=5 OP=0
cfg[2013] = { 1'b0, 8'h67, 8'hb9}; // CH=3 OP=1
cfg[2014] = { 1'b0, 8'h45, 8'h39}; // CH=1 OP=1
cfg[2015] = { 1'b0, 8'h78, 8'he0}; // CH=0 OP=2
cfg[2016] = { 1'b1, 8'hd0, 8'h47}; // CH=3 OP=0
cfg[2017] = { 1'b0, 8'h8b, 8'h89}; // CH=3 OP=2
cfg[2018] = { 1'b1, 8'h9b, 8'h45}; // CH=6 OP=2
cfg[2019] = { 1'b0, 8'hc5, 8'h9f}; // CH=1 OP=1
cfg[2020] = { 1'b0, 8'h4c, 8'hc9}; // CH=0 OP=3
cfg[2021] = { 1'b0, 8'h74, 8'h78}; // CH=0 OP=1
cfg[2022] = { 1'b0, 8'h6e, 8'h70}; // CH=2 OP=3
cfg[2023] = { 1'b1, 8'h62, 8'hd7}; // CH=5 OP=0
cfg[2024] = { 1'b0, 8'ha6, 8'h1d}; // CH=2 OP=1
cfg[2025] = { 1'b1, 8'ha2, 8'h43}; // CH=5 OP=0
cfg[2026] = { 1'b0, 8'h82, 8'hee}; // CH=2 OP=0
cfg[2027] = { 1'b1, 8'hed, 8'h7a}; // CH=4 OP=3
cfg[2028] = { 1'b0, 8'h73, 8'h15}; // CH=3 OP=0
cfg[2029] = { 1'b1, 8'hc0, 8'hda}; // CH=3 OP=0
cfg[2030] = { 1'b0, 8'h38, 8'h54}; // CH=0 OP=2
cfg[2031] = { 1'b1, 8'hb0, 8'hc8}; // CH=3 OP=0
cfg[2032] = { 1'b1, 8'he2, 8'h36}; // CH=5 OP=0
cfg[2033] = { 1'b1, 8'h4c, 8'h98}; // CH=3 OP=3
cfg[2034] = { 1'b0, 8'h97, 8'h3e}; // CH=3 OP=1
cfg[2035] = { 1'b1, 8'h39, 8'h5d}; // CH=4 OP=2
cfg[2036] = { 1'b1, 8'hbc, 8'h4b}; // CH=3 OP=3
cfg[2037] = { 1'b0, 8'ha9, 8'hc5}; // CH=1 OP=2
cfg[2038] = { 1'b0, 8'hd9, 8'hda}; // CH=1 OP=2
cfg[2039] = { 1'b0, 8'h99, 8'h1d}; // CH=1 OP=2
cfg[2040] = { 1'b1, 8'hd1, 8'h71}; // CH=4 OP=0
cfg[2041] = { 1'b0, 8'h82, 8'h3a}; // CH=2 OP=0
cfg[2042] = { 1'b1, 8'h64, 8'h70}; // CH=3 OP=1
cfg[2043] = { 1'b0, 8'hb0, 8'h9}; // CH=0 OP=0
cfg[2044] = { 1'b0, 8'h48, 8'h47}; // CH=0 OP=2
cfg[2045] = { 1'b1, 8'h81, 8'ha4}; // CH=4 OP=0
cfg[2046] = { 1'b0, 8'h3d, 8'hf0}; // CH=1 OP=3
cfg[2047] = { 1'b0, 8'he7, 8'hb5}; // CH=3 OP=1
cfg[2048] = { 1'b0, 8'hb5, 8'h90}; // CH=1 OP=1
cfg[2049] = { 1'b0, 8'h4e, 8'h21}; // CH=2 OP=3
cfg[2050] = { 1'b1, 8'h3f, 8'h92}; // CH=6 OP=3
cfg[2051] = { 1'b0, 8'h3d, 8'ha2}; // CH=1 OP=3
cfg[2052] = { 1'b0, 8'h46, 8'h77}; // CH=2 OP=1
cfg[2053] = { 1'b0, 8'h8d, 8'h84}; // CH=1 OP=3
cfg[2054] = { 1'b0, 8'h32, 8'h7d}; // CH=2 OP=0
cfg[2055] = { 1'b0, 8'hbd, 8'hee}; // CH=1 OP=3
cfg[2056] = { 1'b0, 8'ha4, 8'hd7}; // CH=0 OP=1
cfg[2057] = { 1'b1, 8'ha8, 8'h67}; // CH=3 OP=2
cfg[2058] = { 1'b0, 8'hc9, 8'hac}; // CH=1 OP=2
cfg[2059] = { 1'b1, 8'h5c, 8'hcb}; // CH=3 OP=3
cfg[2060] = { 1'b1, 8'h8b, 8'hb}; // CH=6 OP=2
cfg[2061] = { 1'b0, 8'h91, 8'h65}; // CH=1 OP=0
cfg[2062] = { 1'b1, 8'h47, 8'hab}; // CH=6 OP=1
cfg[2063] = { 1'b1, 8'h46, 8'h39}; // CH=5 OP=1
cfg[2064] = { 1'b1, 8'hc6, 8'h6b}; // CH=5 OP=1
cfg[2065] = { 1'b1, 8'h83, 8'h8d}; // CH=6 OP=0
cfg[2066] = { 1'b1, 8'h34, 8'h64}; // CH=3 OP=1
cfg[2067] = { 1'b0, 8'haf, 8'hd0}; // CH=3 OP=3
cfg[2068] = { 1'b0, 8'h78, 8'h9a}; // CH=0 OP=2
cfg[2069] = { 1'b1, 8'h61, 8'hf6}; // CH=4 OP=0
cfg[2070] = { 1'b0, 8'hec, 8'h1e}; // CH=0 OP=3
cfg[2071] = { 1'b0, 8'h7d, 8'h84}; // CH=1 OP=3
cfg[2072] = { 1'b0, 8'hc4, 8'h2f}; // CH=0 OP=1
cfg[2073] = { 1'b1, 8'hba, 8'h68}; // CH=5 OP=2
cfg[2074] = { 1'b1, 8'h41, 8'hd0}; // CH=4 OP=0
cfg[2075] = { 1'b0, 8'hb1, 8'h54}; // CH=1 OP=0
cfg[2076] = { 1'b1, 8'he5, 8'h7c}; // CH=4 OP=1
cfg[2077] = { 1'b1, 8'h94, 8'h4c}; // CH=3 OP=1
cfg[2078] = { 1'b1, 8'h4c, 8'he6}; // CH=3 OP=3
cfg[2079] = { 1'b0, 8'h9b, 8'h6d}; // CH=3 OP=2
cfg[2080] = { 1'b1, 8'h7f, 8'h59}; // CH=6 OP=3
cfg[2081] = { 1'b0, 8'hae, 8'hf}; // CH=2 OP=3
cfg[2082] = { 1'b1, 8'ha5, 8'h31}; // CH=4 OP=1
cfg[2083] = { 1'b1, 8'h76, 8'hea}; // CH=5 OP=1
cfg[2084] = { 1'b1, 8'hca, 8'h4b}; // CH=5 OP=2
cfg[2085] = { 1'b0, 8'h46, 8'h10}; // CH=2 OP=1
cfg[2086] = { 1'b1, 8'h92, 8'ha1}; // CH=5 OP=0
cfg[2087] = { 1'b0, 8'h79, 8'haa}; // CH=1 OP=2
cfg[2088] = { 1'b0, 8'h55, 8'hf6}; // CH=1 OP=1
cfg[2089] = { 1'b0, 8'h50, 8'h91}; // CH=0 OP=0
cfg[2090] = { 1'b1, 8'hcf, 8'h9b}; // CH=6 OP=3
cfg[2091] = { 1'b0, 8'h7e, 8'haa}; // CH=2 OP=3
cfg[2092] = { 1'b1, 8'h95, 8'hdb}; // CH=4 OP=1
cfg[2093] = { 1'b0, 8'h7f, 8'hc7}; // CH=3 OP=3
cfg[2094] = { 1'b0, 8'hca, 8'hf4}; // CH=2 OP=2
cfg[2095] = { 1'b0, 8'hda, 8'hd2}; // CH=2 OP=2
cfg[2096] = { 1'b0, 8'h7b, 8'h95}; // CH=3 OP=2
cfg[2097] = { 1'b1, 8'hd4, 8'hed}; // CH=3 OP=1
cfg[2098] = { 1'b0, 8'had, 8'h1c}; // CH=1 OP=3
cfg[2099] = { 1'b0, 8'h48, 8'h4f}; // CH=0 OP=2
cfg[2100] = { 1'b1, 8'hf3, 8'h51}; // CH=6 OP=0
cfg[2101] = { 1'b1, 8'hce, 8'hee}; // CH=5 OP=3
cfg[2102] = { 1'b0, 8'h95, 8'h31}; // CH=1 OP=1
cfg[2103] = { 1'b0, 8'h89, 8'he9}; // CH=1 OP=2
cfg[2104] = { 1'b0, 8'h5b, 8'h6c}; // CH=3 OP=2
cfg[2105] = { 1'b1, 8'hf1, 8'h34}; // CH=4 OP=0
cfg[2106] = { 1'b0, 8'hde, 8'h8f}; // CH=2 OP=3
cfg[2107] = { 1'b0, 8'h30, 8'h63}; // CH=0 OP=0
cfg[2108] = { 1'b0, 8'h54, 8'h8d}; // CH=0 OP=1
cfg[2109] = { 1'b1, 8'ha4, 8'h7}; // CH=3 OP=1
cfg[2110] = { 1'b0, 8'hf5, 8'h50}; // CH=1 OP=1
cfg[2111] = { 1'b1, 8'he4, 8'h18}; // CH=3 OP=1
cfg[2112] = { 1'b1, 8'h8b, 8'h74}; // CH=6 OP=2
cfg[2113] = { 1'b0, 8'hf7, 8'hfe}; // CH=3 OP=1
cfg[2114] = { 1'b0, 8'h78, 8'h70}; // CH=0 OP=2
cfg[2115] = { 1'b1, 8'h74, 8'h61}; // CH=3 OP=1
cfg[2116] = { 1'b0, 8'h96, 8'h3f}; // CH=2 OP=1
cfg[2117] = { 1'b0, 8'hd4, 8'h70}; // CH=0 OP=1
cfg[2118] = { 1'b1, 8'hc0, 8'hc4}; // CH=3 OP=0
cfg[2119] = { 1'b0, 8'hf4, 8'h68}; // CH=0 OP=1
cfg[2120] = { 1'b0, 8'h8e, 8'h5e}; // CH=2 OP=3
cfg[2121] = { 1'b0, 8'h57, 8'h10}; // CH=3 OP=1
cfg[2122] = { 1'b1, 8'h55, 8'h53}; // CH=4 OP=1
cfg[2123] = { 1'b0, 8'hc0, 8'h4a}; // CH=0 OP=0
cfg[2124] = { 1'b0, 8'h5f, 8'hc2}; // CH=3 OP=3
cfg[2125] = { 1'b1, 8'h8d, 8'h37}; // CH=4 OP=3
cfg[2126] = { 1'b0, 8'h30, 8'hcd}; // CH=0 OP=0
cfg[2127] = { 1'b0, 8'hf5, 8'h3e}; // CH=1 OP=1
cfg[2128] = { 1'b0, 8'h5d, 8'h64}; // CH=1 OP=3
cfg[2129] = { 1'b0, 8'hbb, 8'hdb}; // CH=3 OP=2
cfg[2130] = { 1'b1, 8'hfd, 8'h69}; // CH=4 OP=3
cfg[2131] = { 1'b1, 8'h54, 8'h6c}; // CH=3 OP=1
cfg[2132] = { 1'b1, 8'haa, 8'hc0}; // CH=5 OP=2
cfg[2133] = { 1'b1, 8'h6a, 8'ha}; // CH=5 OP=2
cfg[2134] = { 1'b1, 8'hc9, 8'hcd}; // CH=4 OP=2
cfg[2135] = { 1'b0, 8'h56, 8'h4}; // CH=2 OP=1
cfg[2136] = { 1'b0, 8'h76, 8'hd1}; // CH=2 OP=1
cfg[2137] = { 1'b1, 8'hb4, 8'h73}; // CH=3 OP=1
cfg[2138] = { 1'b0, 8'hb1, 8'hd5}; // CH=1 OP=0
cfg[2139] = { 1'b1, 8'h6d, 8'hf4}; // CH=4 OP=3
cfg[2140] = { 1'b0, 8'h6a, 8'h5d}; // CH=2 OP=2
cfg[2141] = { 1'b0, 8'hbf, 8'hca}; // CH=3 OP=3
cfg[2142] = { 1'b1, 8'h69, 8'h8a}; // CH=4 OP=2
cfg[2143] = { 1'b0, 8'hd3, 8'h94}; // CH=3 OP=0
cfg[2144] = { 1'b1, 8'h9c, 8'h61}; // CH=3 OP=3
cfg[2145] = { 1'b1, 8'hf2, 8'h65}; // CH=5 OP=0
cfg[2146] = { 1'b1, 8'h68, 8'h37}; // CH=3 OP=2
cfg[2147] = { 1'b0, 8'h44, 8'haa}; // CH=0 OP=1
cfg[2148] = { 1'b0, 8'hf6, 8'h36}; // CH=2 OP=1
cfg[2149] = { 1'b1, 8'h63, 8'h2a}; // CH=6 OP=0
cfg[2150] = { 1'b0, 8'hcd, 8'h87}; // CH=1 OP=3
cfg[2151] = { 1'b0, 8'h8c, 8'h51}; // CH=0 OP=3
cfg[2152] = { 1'b1, 8'hf5, 8'hdb}; // CH=4 OP=1
cfg[2153] = { 1'b1, 8'hc8, 8'h70}; // CH=3 OP=2
cfg[2154] = { 1'b0, 8'h64, 8'hd1}; // CH=0 OP=1
cfg[2155] = { 1'b1, 8'h57, 8'h37}; // CH=6 OP=1
cfg[2156] = { 1'b0, 8'hbf, 8'h6e}; // CH=3 OP=3
cfg[2157] = { 1'b1, 8'hdc, 8'h18}; // CH=3 OP=3
cfg[2158] = { 1'b1, 8'hbd, 8'h98}; // CH=4 OP=3
cfg[2159] = { 1'b0, 8'h8c, 8'h3c}; // CH=0 OP=3
cfg[2160] = { 1'b0, 8'hf2, 8'hee}; // CH=2 OP=0
cfg[2161] = { 1'b1, 8'h93, 8'h7a}; // CH=6 OP=0
cfg[2162] = { 1'b1, 8'h3c, 8'h70}; // CH=3 OP=3
cfg[2163] = { 1'b1, 8'hda, 8'h38}; // CH=5 OP=2
cfg[2164] = { 1'b0, 8'hdb, 8'h9d}; // CH=3 OP=2
cfg[2165] = { 1'b1, 8'h6d, 8'hf4}; // CH=4 OP=3
cfg[2166] = { 1'b1, 8'hf0, 8'hb3}; // CH=3 OP=0
cfg[2167] = { 1'b0, 8'hb8, 8'h90}; // CH=0 OP=2
cfg[2168] = { 1'b0, 8'h75, 8'ha2}; // CH=1 OP=1
cfg[2169] = { 1'b0, 8'h96, 8'hdf}; // CH=2 OP=1
cfg[2170] = { 1'b0, 8'h84, 8'ha3}; // CH=0 OP=1
cfg[2171] = { 1'b0, 8'hfe, 8'hb8}; // CH=2 OP=3
cfg[2172] = { 1'b1, 8'h6e, 8'ha9}; // CH=5 OP=3
cfg[2173] = { 1'b1, 8'ha7, 8'ha}; // CH=6 OP=1
cfg[2174] = { 1'b1, 8'h44, 8'h3d}; // CH=3 OP=1
cfg[2175] = { 1'b0, 8'h38, 8'ha6}; // CH=0 OP=2
cfg[2176] = { 1'b0, 8'heb, 8'h7e}; // CH=3 OP=2
cfg[2177] = { 1'b0, 8'h7b, 8'h6e}; // CH=3 OP=2
cfg[2178] = { 1'b0, 8'h5a, 8'hf6}; // CH=2 OP=2
cfg[2179] = { 1'b1, 8'hf0, 8'hfd}; // CH=3 OP=0
cfg[2180] = { 1'b1, 8'h74, 8'ha0}; // CH=3 OP=1
cfg[2181] = { 1'b0, 8'h72, 8'h58}; // CH=2 OP=0
cfg[2182] = { 1'b1, 8'he1, 8'h2}; // CH=4 OP=0
cfg[2183] = { 1'b1, 8'h88, 8'hc}; // CH=3 OP=2
cfg[2184] = { 1'b0, 8'hcc, 8'h49}; // CH=0 OP=3
cfg[2185] = { 1'b1, 8'h5b, 8'hf0}; // CH=6 OP=2
cfg[2186] = { 1'b0, 8'h87, 8'hef}; // CH=3 OP=1
cfg[2187] = { 1'b0, 8'h6c, 8'h6b}; // CH=0 OP=3
cfg[2188] = { 1'b0, 8'hc6, 8'h89}; // CH=2 OP=1
cfg[2189] = { 1'b1, 8'hb6, 8'h86}; // CH=5 OP=1
cfg[2190] = { 1'b1, 8'h7e, 8'h26}; // CH=5 OP=3
cfg[2191] = { 1'b0, 8'h80, 8'h5a}; // CH=0 OP=0
cfg[2192] = { 1'b1, 8'h8d, 8'hb7}; // CH=4 OP=3
cfg[2193] = { 1'b1, 8'hd6, 8'h8}; // CH=5 OP=1
cfg[2194] = { 1'b1, 8'hc6, 8'h27}; // CH=5 OP=1
cfg[2195] = { 1'b1, 8'h34, 8'h82}; // CH=3 OP=1
cfg[2196] = { 1'b1, 8'h30, 8'h9}; // CH=3 OP=0
cfg[2197] = { 1'b1, 8'hb9, 8'he3}; // CH=4 OP=2
cfg[2198] = { 1'b1, 8'h3f, 8'h78}; // CH=6 OP=3
cfg[2199] = { 1'b1, 8'h65, 8'h29}; // CH=4 OP=1
cfg[2200] = { 1'b1, 8'he3, 8'h40}; // CH=6 OP=0
cfg[2201] = { 1'b0, 8'h64, 8'h9b}; // CH=0 OP=1
cfg[2202] = { 1'b1, 8'hf1, 8'h52}; // CH=4 OP=0
cfg[2203] = { 1'b1, 8'hc7, 8'h5a}; // CH=6 OP=1
cfg[2204] = { 1'b0, 8'h8e, 8'h81}; // CH=2 OP=3
cfg[2205] = { 1'b0, 8'hc2, 8'h3}; // CH=2 OP=0
cfg[2206] = { 1'b1, 8'hd3, 8'hd}; // CH=6 OP=0
cfg[2207] = { 1'b1, 8'hb6, 8'h82}; // CH=5 OP=1
cfg[2208] = { 1'b0, 8'hcf, 8'hbe}; // CH=3 OP=3
cfg[2209] = { 1'b1, 8'h34, 8'h58}; // CH=3 OP=1
cfg[2210] = { 1'b1, 8'h83, 8'h98}; // CH=6 OP=0
cfg[2211] = { 1'b1, 8'hb8, 8'h7b}; // CH=3 OP=2
cfg[2212] = { 1'b0, 8'hf3, 8'h6c}; // CH=3 OP=0
cfg[2213] = { 1'b0, 8'h62, 8'h34}; // CH=2 OP=0
cfg[2214] = { 1'b0, 8'h65, 8'he2}; // CH=1 OP=1
cfg[2215] = { 1'b0, 8'h72, 8'h89}; // CH=2 OP=0
cfg[2216] = { 1'b1, 8'hf5, 8'h60}; // CH=4 OP=1
cfg[2217] = { 1'b1, 8'hb3, 8'hf0}; // CH=6 OP=0
cfg[2218] = { 1'b0, 8'h62, 8'hbf}; // CH=2 OP=0
cfg[2219] = { 1'b0, 8'hb0, 8'hf3}; // CH=0 OP=0
cfg[2220] = { 1'b0, 8'h69, 8'h86}; // CH=1 OP=2
cfg[2221] = { 1'b0, 8'h5c, 8'hf2}; // CH=0 OP=3
cfg[2222] = { 1'b0, 8'h5c, 8'h26}; // CH=0 OP=3
cfg[2223] = { 1'b0, 8'h3e, 8'he8}; // CH=2 OP=3
cfg[2224] = { 1'b0, 8'hc7, 8'h6d}; // CH=3 OP=1
cfg[2225] = { 1'b0, 8'hf5, 8'hc4}; // CH=1 OP=1
cfg[2226] = { 1'b0, 8'ha8, 8'h17}; // CH=0 OP=2
cfg[2227] = { 1'b0, 8'ha2, 8'hd6}; // CH=2 OP=0
cfg[2228] = { 1'b1, 8'hce, 8'h38}; // CH=5 OP=3
cfg[2229] = { 1'b0, 8'h5a, 8'he9}; // CH=2 OP=2
cfg[2230] = { 1'b0, 8'h4c, 8'h14}; // CH=0 OP=3
cfg[2231] = { 1'b0, 8'h73, 8'hdb}; // CH=3 OP=0
cfg[2232] = { 1'b1, 8'h5b, 8'h3}; // CH=6 OP=2
cfg[2233] = { 1'b1, 8'hc8, 8'h91}; // CH=3 OP=2
cfg[2234] = { 1'b1, 8'h8d, 8'h92}; // CH=4 OP=3
cfg[2235] = { 1'b0, 8'h5f, 8'h87}; // CH=3 OP=3
cfg[2236] = { 1'b0, 8'h6d, 8'h30}; // CH=1 OP=3
cfg[2237] = { 1'b0, 8'hf0, 8'h3b}; // CH=0 OP=0
cfg[2238] = { 1'b1, 8'hc4, 8'hdd}; // CH=3 OP=1
cfg[2239] = { 1'b0, 8'hae, 8'hc}; // CH=2 OP=3
cfg[2240] = { 1'b0, 8'h5d, 8'h6a}; // CH=1 OP=3
cfg[2241] = { 1'b1, 8'h68, 8'hdd}; // CH=3 OP=2
cfg[2242] = { 1'b1, 8'hb1, 8'h39}; // CH=4 OP=0
cfg[2243] = { 1'b0, 8'hc2, 8'h1}; // CH=2 OP=0
cfg[2244] = { 1'b0, 8'hfb, 8'h8e}; // CH=3 OP=2
cfg[2245] = { 1'b0, 8'h4b, 8'hed}; // CH=3 OP=2
cfg[2246] = { 1'b0, 8'h71, 8'h5a}; // CH=1 OP=0
cfg[2247] = { 1'b1, 8'h61, 8'h69}; // CH=4 OP=0
cfg[2248] = { 1'b0, 8'he5, 8'h47}; // CH=1 OP=1
cfg[2249] = { 1'b1, 8'h93, 8'h43}; // CH=6 OP=0
cfg[2250] = { 1'b1, 8'hf0, 8'hae}; // CH=3 OP=0
cfg[2251] = { 1'b1, 8'h58, 8'h8b}; // CH=3 OP=2
cfg[2252] = { 1'b0, 8'hfe, 8'hc4}; // CH=2 OP=3
cfg[2253] = { 1'b0, 8'h54, 8'hcc}; // CH=0 OP=1
cfg[2254] = { 1'b1, 8'h42, 8'hcb}; // CH=5 OP=0
cfg[2255] = { 1'b0, 8'h9c, 8'ha5}; // CH=0 OP=3
cfg[2256] = { 1'b0, 8'he5, 8'hba}; // CH=1 OP=1
cfg[2257] = { 1'b0, 8'ha0, 8'h4d}; // CH=0 OP=0
cfg[2258] = { 1'b0, 8'hfc, 8'hbb}; // CH=0 OP=3
cfg[2259] = { 1'b1, 8'h88, 8'h82}; // CH=3 OP=2
cfg[2260] = { 1'b0, 8'h4c, 8'hf0}; // CH=0 OP=3
cfg[2261] = { 1'b0, 8'hda, 8'hef}; // CH=2 OP=2
cfg[2262] = { 1'b0, 8'ha2, 8'h67}; // CH=2 OP=0
cfg[2263] = { 1'b1, 8'hb4, 8'ha9}; // CH=3 OP=1
cfg[2264] = { 1'b0, 8'h38, 8'h45}; // CH=0 OP=2
cfg[2265] = { 1'b0, 8'h7c, 8'h4b}; // CH=0 OP=3
cfg[2266] = { 1'b0, 8'ha4, 8'h29}; // CH=0 OP=1
cfg[2267] = { 1'b0, 8'h5f, 8'h77}; // CH=3 OP=3
cfg[2268] = { 1'b0, 8'hce, 8'h74}; // CH=2 OP=3
cfg[2269] = { 1'b0, 8'hbf, 8'he}; // CH=3 OP=3
cfg[2270] = { 1'b0, 8'hae, 8'h1c}; // CH=2 OP=3
cfg[2271] = { 1'b1, 8'hbe, 8'hf7}; // CH=5 OP=3
cfg[2272] = { 1'b0, 8'h99, 8'h99}; // CH=1 OP=2
cfg[2273] = { 1'b1, 8'hb0, 8'h4d}; // CH=3 OP=0
cfg[2274] = { 1'b0, 8'hfc, 8'h53}; // CH=0 OP=3
cfg[2275] = { 1'b0, 8'h94, 8'hcf}; // CH=0 OP=1
cfg[2276] = { 1'b1, 8'hcd, 8'h73}; // CH=4 OP=3
cfg[2277] = { 1'b0, 8'hb8, 8'hd2}; // CH=0 OP=2
cfg[2278] = { 1'b1, 8'hb4, 8'he7}; // CH=3 OP=1
cfg[2279] = { 1'b1, 8'hfd, 8'ha6}; // CH=4 OP=3
cfg[2280] = { 1'b0, 8'h58, 8'h54}; // CH=0 OP=2
cfg[2281] = { 1'b1, 8'h98, 8'h12}; // CH=3 OP=2
cfg[2282] = { 1'b1, 8'he5, 8'h85}; // CH=4 OP=1
cfg[2283] = { 1'b0, 8'h6b, 8'h35}; // CH=3 OP=2
cfg[2284] = { 1'b1, 8'he7, 8'h31}; // CH=6 OP=1
cfg[2285] = { 1'b0, 8'h5a, 8'hdc}; // CH=2 OP=2
cfg[2286] = { 1'b1, 8'hac, 8'h21}; // CH=3 OP=3
cfg[2287] = { 1'b1, 8'h93, 8'ha}; // CH=6 OP=0
cfg[2288] = { 1'b0, 8'h3a, 8'hf5}; // CH=2 OP=2
cfg[2289] = { 1'b1, 8'h8e, 8'hfd}; // CH=5 OP=3
cfg[2290] = { 1'b1, 8'ha1, 8'hfc}; // CH=4 OP=0
cfg[2291] = { 1'b1, 8'h4c, 8'h94}; // CH=3 OP=3
cfg[2292] = { 1'b0, 8'hb7, 8'h7a}; // CH=3 OP=1
cfg[2293] = { 1'b1, 8'he9, 8'h28}; // CH=4 OP=2
cfg[2294] = { 1'b1, 8'haf, 8'hf}; // CH=6 OP=3
cfg[2295] = { 1'b1, 8'h42, 8'h6a}; // CH=5 OP=0
cfg[2296] = { 1'b0, 8'hee, 8'h97}; // CH=2 OP=3
cfg[2297] = { 1'b0, 8'h81, 8'ha1}; // CH=1 OP=0
cfg[2298] = { 1'b0, 8'hbb, 8'h96}; // CH=3 OP=2
cfg[2299] = { 1'b1, 8'h4a, 8'h94}; // CH=5 OP=2
cfg[2300] = { 1'b0, 8'heb, 8'h90}; // CH=3 OP=2
cfg[2301] = { 1'b1, 8'h37, 8'h25}; // CH=6 OP=1
cfg[2302] = { 1'b1, 8'h48, 8'h9f}; // CH=3 OP=2
cfg[2303] = { 1'b0, 8'h71, 8'h84}; // CH=1 OP=0
cfg[2304] = { 1'b1, 8'h80, 8'h79}; // CH=3 OP=0
cfg[2305] = { 1'b0, 8'hea, 8'h4b}; // CH=2 OP=2
cfg[2306] = { 1'b0, 8'h81, 8'h3d}; // CH=1 OP=0
cfg[2307] = { 1'b0, 8'h48, 8'h9}; // CH=0 OP=2
cfg[2308] = { 1'b1, 8'h48, 8'hb9}; // CH=3 OP=2
cfg[2309] = { 1'b1, 8'hdd, 8'h4d}; // CH=4 OP=3
cfg[2310] = { 1'b0, 8'h70, 8'hd5}; // CH=0 OP=0
cfg[2311] = { 1'b0, 8'hb8, 8'ha1}; // CH=0 OP=2
cfg[2312] = { 1'b1, 8'h9f, 8'h26}; // CH=6 OP=3
cfg[2313] = { 1'b0, 8'hea, 8'h99}; // CH=2 OP=2
cfg[2314] = { 1'b0, 8'h38, 8'h71}; // CH=0 OP=2
cfg[2315] = { 1'b1, 8'h80, 8'h38}; // CH=3 OP=0
cfg[2316] = { 1'b1, 8'h83, 8'hf1}; // CH=6 OP=0
cfg[2317] = { 1'b1, 8'hd1, 8'h3e}; // CH=4 OP=0
cfg[2318] = { 1'b0, 8'hc3, 8'h1c}; // CH=3 OP=0
cfg[2319] = { 1'b0, 8'he0, 8'h79}; // CH=0 OP=0
cfg[2320] = { 1'b0, 8'hfb, 8'h32}; // CH=3 OP=2
cfg[2321] = { 1'b0, 8'hfd, 8'h5b}; // CH=1 OP=3
cfg[2322] = { 1'b1, 8'h96, 8'h5}; // CH=5 OP=1
cfg[2323] = { 1'b0, 8'h98, 8'h9a}; // CH=0 OP=2
cfg[2324] = { 1'b0, 8'hc9, 8'h40}; // CH=1 OP=2
cfg[2325] = { 1'b0, 8'h5e, 8'hc0}; // CH=2 OP=3
cfg[2326] = { 1'b0, 8'h3c, 8'h43}; // CH=0 OP=3
cfg[2327] = { 1'b0, 8'h34, 8'h14}; // CH=0 OP=1
cfg[2328] = { 1'b0, 8'h53, 8'hed}; // CH=3 OP=0
cfg[2329] = { 1'b1, 8'hc9, 8'hcd}; // CH=4 OP=2
cfg[2330] = { 1'b0, 8'hc6, 8'hf9}; // CH=2 OP=1
cfg[2331] = { 1'b0, 8'h5c, 8'h2a}; // CH=0 OP=3
cfg[2332] = { 1'b0, 8'h64, 8'hc4}; // CH=0 OP=1
cfg[2333] = { 1'b0, 8'ha4, 8'h74}; // CH=0 OP=1
cfg[2334] = { 1'b0, 8'h64, 8'h5d}; // CH=0 OP=1
cfg[2335] = { 1'b0, 8'ha8, 8'h37}; // CH=0 OP=2
cfg[2336] = { 1'b0, 8'hbc, 8'h4f}; // CH=0 OP=3
cfg[2337] = { 1'b0, 8'hda, 8'h84}; // CH=2 OP=2
cfg[2338] = { 1'b0, 8'h72, 8'hd7}; // CH=2 OP=0
cfg[2339] = { 1'b1, 8'h3b, 8'hea}; // CH=6 OP=2
cfg[2340] = { 1'b0, 8'h60, 8'he3}; // CH=0 OP=0
cfg[2341] = { 1'b0, 8'h8b, 8'h61}; // CH=3 OP=2
cfg[2342] = { 1'b0, 8'h4f, 8'h50}; // CH=3 OP=3
cfg[2343] = { 1'b1, 8'hc4, 8'hd6}; // CH=3 OP=1
cfg[2344] = { 1'b1, 8'hd5, 8'h26}; // CH=4 OP=1
cfg[2345] = { 1'b0, 8'hbf, 8'hd0}; // CH=3 OP=3
cfg[2346] = { 1'b1, 8'hd4, 8'h8c}; // CH=3 OP=1
cfg[2347] = { 1'b1, 8'hd6, 8'h67}; // CH=5 OP=1
cfg[2348] = { 1'b0, 8'ha5, 8'hd9}; // CH=1 OP=1
cfg[2349] = { 1'b0, 8'h3d, 8'h14}; // CH=1 OP=3
cfg[2350] = { 1'b1, 8'h9b, 8'h75}; // CH=6 OP=2
cfg[2351] = { 1'b1, 8'h56, 8'h0}; // CH=5 OP=1
cfg[2352] = { 1'b1, 8'h75, 8'h4f}; // CH=4 OP=1
cfg[2353] = { 1'b1, 8'h38, 8'h13}; // CH=3 OP=2
cfg[2354] = { 1'b0, 8'h60, 8'h34}; // CH=0 OP=0
cfg[2355] = { 1'b1, 8'h30, 8'h8c}; // CH=3 OP=0
cfg[2356] = { 1'b0, 8'hbd, 8'h34}; // CH=1 OP=3
cfg[2357] = { 1'b0, 8'hbc, 8'h5f}; // CH=0 OP=3
cfg[2358] = { 1'b0, 8'h62, 8'hfd}; // CH=2 OP=0
cfg[2359] = { 1'b0, 8'h9f, 8'h11}; // CH=3 OP=3
cfg[2360] = { 1'b0, 8'h3b, 8'h86}; // CH=3 OP=2
cfg[2361] = { 1'b1, 8'h91, 8'h86}; // CH=4 OP=0
cfg[2362] = { 1'b0, 8'he9, 8'hd6}; // CH=1 OP=2
cfg[2363] = { 1'b0, 8'h9f, 8'ha5}; // CH=3 OP=3
cfg[2364] = { 1'b0, 8'hcf, 8'haa}; // CH=3 OP=3
cfg[2365] = { 1'b1, 8'h8c, 8'hde}; // CH=3 OP=3
cfg[2366] = { 1'b1, 8'hb0, 8'h3e}; // CH=3 OP=0
cfg[2367] = { 1'b0, 8'had, 8'ha0}; // CH=1 OP=3
cfg[2368] = { 1'b0, 8'hbf, 8'hee}; // CH=3 OP=3
cfg[2369] = { 1'b1, 8'h45, 8'hc}; // CH=4 OP=1
cfg[2370] = { 1'b0, 8'hcc, 8'h5b}; // CH=0 OP=3
cfg[2371] = { 1'b1, 8'ha2, 8'h2b}; // CH=5 OP=0
cfg[2372] = { 1'b1, 8'h8b, 8'h53}; // CH=6 OP=2
cfg[2373] = { 1'b0, 8'ha9, 8'hf8}; // CH=1 OP=2
cfg[2374] = { 1'b1, 8'h54, 8'hf1}; // CH=3 OP=1
cfg[2375] = { 1'b0, 8'h32, 8'hfc}; // CH=2 OP=0
cfg[2376] = { 1'b1, 8'h70, 8'hed}; // CH=3 OP=0
cfg[2377] = { 1'b1, 8'hab, 8'h9b}; // CH=6 OP=2
cfg[2378] = { 1'b1, 8'h5b, 8'hd8}; // CH=6 OP=2
cfg[2379] = { 1'b1, 8'h45, 8'h1d}; // CH=4 OP=1
cfg[2380] = { 1'b1, 8'hc1, 8'he9}; // CH=4 OP=0
cfg[2381] = { 1'b0, 8'h42, 8'h8b}; // CH=2 OP=0
cfg[2382] = { 1'b1, 8'hde, 8'h17}; // CH=5 OP=3
cfg[2383] = { 1'b0, 8'hcf, 8'h61}; // CH=3 OP=3
cfg[2384] = { 1'b0, 8'hcb, 8'h90}; // CH=3 OP=2
cfg[2385] = { 1'b1, 8'hb8, 8'h4b}; // CH=3 OP=2
cfg[2386] = { 1'b1, 8'h54, 8'hb6}; // CH=3 OP=1
cfg[2387] = { 1'b0, 8'hff, 8'hcf}; // CH=3 OP=3
cfg[2388] = { 1'b1, 8'h5a, 8'ha7}; // CH=5 OP=2
cfg[2389] = { 1'b0, 8'ha0, 8'hc5}; // CH=0 OP=0
cfg[2390] = { 1'b1, 8'h61, 8'hae}; // CH=4 OP=0
cfg[2391] = { 1'b0, 8'ha3, 8'h3a}; // CH=3 OP=0
cfg[2392] = { 1'b1, 8'ha6, 8'h51}; // CH=5 OP=1
cfg[2393] = { 1'b1, 8'h5e, 8'h11}; // CH=5 OP=3
cfg[2394] = { 1'b0, 8'h6d, 8'h97}; // CH=1 OP=3
cfg[2395] = { 1'b0, 8'h99, 8'he2}; // CH=1 OP=2
cfg[2396] = { 1'b0, 8'h68, 8'hec}; // CH=0 OP=2
cfg[2397] = { 1'b1, 8'h90, 8'hb3}; // CH=3 OP=0
cfg[2398] = { 1'b0, 8'h30, 8'hd5}; // CH=0 OP=0
cfg[2399] = { 1'b1, 8'h91, 8'h83}; // CH=4 OP=0
cfg[2400] = { 1'b1, 8'h34, 8'hbd}; // CH=3 OP=1
cfg[2401] = { 1'b1, 8'hda, 8'he}; // CH=5 OP=2
cfg[2402] = { 1'b0, 8'he2, 8'h20}; // CH=2 OP=0
cfg[2403] = { 1'b1, 8'h79, 8'h46}; // CH=4 OP=2
cfg[2404] = { 1'b0, 8'h5c, 8'hb3}; // CH=0 OP=3
cfg[2405] = { 1'b0, 8'hf5, 8'hd7}; // CH=1 OP=1
cfg[2406] = { 1'b0, 8'h5d, 8'hc4}; // CH=1 OP=3
cfg[2407] = { 1'b0, 8'h6d, 8'h77}; // CH=1 OP=3
cfg[2408] = { 1'b0, 8'h42, 8'hfd}; // CH=2 OP=0
cfg[2409] = { 1'b0, 8'hc6, 8'hbd}; // CH=2 OP=1
cfg[2410] = { 1'b1, 8'h83, 8'h48}; // CH=6 OP=0
cfg[2411] = { 1'b1, 8'h92, 8'h85}; // CH=5 OP=0
cfg[2412] = { 1'b0, 8'hb2, 8'h52}; // CH=2 OP=0
cfg[2413] = { 1'b0, 8'hf8, 8'h7d}; // CH=0 OP=2
cfg[2414] = { 1'b1, 8'hab, 8'hd1}; // CH=6 OP=2
cfg[2415] = { 1'b1, 8'h82, 8'h8}; // CH=5 OP=0
cfg[2416] = { 1'b0, 8'h46, 8'h74}; // CH=2 OP=1
cfg[2417] = { 1'b0, 8'hbe, 8'h16}; // CH=2 OP=3
cfg[2418] = { 1'b1, 8'hbb, 8'h48}; // CH=6 OP=2
cfg[2419] = { 1'b0, 8'h78, 8'haa}; // CH=0 OP=2
cfg[2420] = { 1'b0, 8'hc1, 8'h9d}; // CH=1 OP=0
cfg[2421] = { 1'b1, 8'h46, 8'hc5}; // CH=5 OP=1
cfg[2422] = { 1'b1, 8'h98, 8'hc7}; // CH=3 OP=2
cfg[2423] = { 1'b1, 8'h41, 8'hab}; // CH=4 OP=0
cfg[2424] = { 1'b0, 8'hec, 8'he7}; // CH=0 OP=3
cfg[2425] = { 1'b0, 8'h6f, 8'hef}; // CH=3 OP=3
cfg[2426] = { 1'b0, 8'hb5, 8'h63}; // CH=1 OP=1
cfg[2427] = { 1'b0, 8'h73, 8'h7a}; // CH=3 OP=0
cfg[2428] = { 1'b0, 8'hb2, 8'hc2}; // CH=2 OP=0
cfg[2429] = { 1'b1, 8'h34, 8'ha7}; // CH=3 OP=1
cfg[2430] = { 1'b0, 8'h39, 8'h68}; // CH=1 OP=2
cfg[2431] = { 1'b1, 8'hd1, 8'haf}; // CH=4 OP=0
cfg[2432] = { 1'b0, 8'h41, 8'h47}; // CH=1 OP=0
cfg[2433] = { 1'b1, 8'h4a, 8'h5c}; // CH=5 OP=2
cfg[2434] = { 1'b0, 8'h33, 8'h48}; // CH=3 OP=0
cfg[2435] = { 1'b1, 8'h96, 8'h7c}; // CH=5 OP=1
cfg[2436] = { 1'b1, 8'he0, 8'hf9}; // CH=3 OP=0
cfg[2437] = { 1'b1, 8'ha1, 8'hd3}; // CH=4 OP=0
cfg[2438] = { 1'b0, 8'hd5, 8'hb7}; // CH=1 OP=1
cfg[2439] = { 1'b0, 8'hce, 8'h1f}; // CH=2 OP=3
cfg[2440] = { 1'b1, 8'hfa, 8'hb0}; // CH=5 OP=2
cfg[2441] = { 1'b0, 8'h56, 8'h73}; // CH=2 OP=1
cfg[2442] = { 1'b0, 8'h9e, 8'hb7}; // CH=2 OP=3
cfg[2443] = { 1'b0, 8'h56, 8'hea}; // CH=2 OP=1
cfg[2444] = { 1'b0, 8'hc3, 8'h80}; // CH=3 OP=0
cfg[2445] = { 1'b1, 8'ha3, 8'h91}; // CH=6 OP=0
cfg[2446] = { 1'b0, 8'hb3, 8'h64}; // CH=3 OP=0
cfg[2447] = { 1'b1, 8'h6a, 8'ha4}; // CH=5 OP=2
cfg[2448] = { 1'b0, 8'h89, 8'hee}; // CH=1 OP=2
cfg[2449] = { 1'b1, 8'h58, 8'h8}; // CH=3 OP=2
cfg[2450] = { 1'b0, 8'h6e, 8'hb9}; // CH=2 OP=3
cfg[2451] = { 1'b0, 8'he1, 8'hab}; // CH=1 OP=0
cfg[2452] = { 1'b0, 8'h98, 8'he7}; // CH=0 OP=2
cfg[2453] = { 1'b1, 8'h82, 8'h2f}; // CH=5 OP=0
cfg[2454] = { 1'b1, 8'hb1, 8'hf3}; // CH=4 OP=0
cfg[2455] = { 1'b1, 8'h5d, 8'hbb}; // CH=4 OP=3
cfg[2456] = { 1'b1, 8'hab, 8'h6e}; // CH=6 OP=2
cfg[2457] = { 1'b1, 8'hcd, 8'hd8}; // CH=4 OP=3
cfg[2458] = { 1'b0, 8'hfe, 8'h62}; // CH=2 OP=3
cfg[2459] = { 1'b0, 8'h4b, 8'hba}; // CH=3 OP=2
cfg[2460] = { 1'b0, 8'hf6, 8'h19}; // CH=2 OP=1
cfg[2461] = { 1'b1, 8'hdd, 8'h7a}; // CH=4 OP=3
cfg[2462] = { 1'b1, 8'hce, 8'h79}; // CH=5 OP=3
cfg[2463] = { 1'b0, 8'he6, 8'h25}; // CH=2 OP=1
cfg[2464] = { 1'b1, 8'ha1, 8'hb9}; // CH=4 OP=0
cfg[2465] = { 1'b0, 8'hb9, 8'hb0}; // CH=1 OP=2
cfg[2466] = { 1'b0, 8'h87, 8'he8}; // CH=3 OP=1
cfg[2467] = { 1'b0, 8'h85, 8'h4a}; // CH=1 OP=1
cfg[2468] = { 1'b0, 8'h94, 8'h4}; // CH=0 OP=1
cfg[2469] = { 1'b0, 8'hae, 8'h2c}; // CH=2 OP=3
cfg[2470] = { 1'b0, 8'h88, 8'h35}; // CH=0 OP=2
cfg[2471] = { 1'b0, 8'h94, 8'ha1}; // CH=0 OP=1
cfg[2472] = { 1'b1, 8'h94, 8'h6f}; // CH=3 OP=1
cfg[2473] = { 1'b1, 8'h45, 8'h55}; // CH=4 OP=1
cfg[2474] = { 1'b0, 8'h54, 8'hf6}; // CH=0 OP=1
cfg[2475] = { 1'b0, 8'hd4, 8'h6}; // CH=0 OP=1
cfg[2476] = { 1'b1, 8'haa, 8'h94}; // CH=5 OP=2
cfg[2477] = { 1'b1, 8'h3e, 8'h1a}; // CH=5 OP=3
cfg[2478] = { 1'b0, 8'h6a, 8'hc7}; // CH=2 OP=2
cfg[2479] = { 1'b0, 8'ha0, 8'h71}; // CH=0 OP=0
cfg[2480] = { 1'b0, 8'h76, 8'hf9}; // CH=2 OP=1
cfg[2481] = { 1'b1, 8'h70, 8'h8e}; // CH=3 OP=0
cfg[2482] = { 1'b0, 8'h8f, 8'h22}; // CH=3 OP=3
cfg[2483] = { 1'b1, 8'h67, 8'h68}; // CH=6 OP=1
cfg[2484] = { 1'b0, 8'hef, 8'hbc}; // CH=3 OP=3
cfg[2485] = { 1'b0, 8'hc4, 8'hc9}; // CH=0 OP=1
cfg[2486] = { 1'b1, 8'h6e, 8'h5e}; // CH=5 OP=3
cfg[2487] = { 1'b1, 8'h81, 8'h78}; // CH=4 OP=0
cfg[2488] = { 1'b1, 8'h48, 8'h26}; // CH=3 OP=2
cfg[2489] = { 1'b1, 8'hba, 8'h83}; // CH=5 OP=2
cfg[2490] = { 1'b1, 8'hb3, 8'h7}; // CH=6 OP=0
cfg[2491] = { 1'b0, 8'h41, 8'h2d}; // CH=1 OP=0
cfg[2492] = { 1'b0, 8'h64, 8'hc1}; // CH=0 OP=1
cfg[2493] = { 1'b1, 8'hcc, 8'hab}; // CH=3 OP=3
cfg[2494] = { 1'b0, 8'h88, 8'h8b}; // CH=0 OP=2
cfg[2495] = { 1'b1, 8'h51, 8'h71}; // CH=4 OP=0
cfg[2496] = { 1'b1, 8'haf, 8'h47}; // CH=6 OP=3
cfg[2497] = { 1'b0, 8'hd7, 8'h56}; // CH=3 OP=1
cfg[2498] = { 1'b1, 8'h5a, 8'h4e}; // CH=5 OP=2
cfg[2499] = { 1'b1, 8'hb2, 8'hda}; // CH=5 OP=0
cfg[2500] = { 1'b0, 8'h80, 8'h8d}; // CH=0 OP=0
cfg[2501] = { 1'b1, 8'hbe, 8'hcf}; // CH=5 OP=3
cfg[2502] = { 1'b1, 8'h8b, 8'h33}; // CH=6 OP=2
cfg[2503] = { 1'b0, 8'hbf, 8'hff}; // CH=3 OP=3
cfg[2504] = { 1'b1, 8'he2, 8'h87}; // CH=5 OP=0
cfg[2505] = { 1'b0, 8'hca, 8'hd8}; // CH=2 OP=2
cfg[2506] = { 1'b1, 8'haf, 8'h88}; // CH=6 OP=3
cfg[2507] = { 1'b1, 8'hfd, 8'hae}; // CH=4 OP=3
cfg[2508] = { 1'b1, 8'hce, 8'h9}; // CH=5 OP=3
cfg[2509] = { 1'b1, 8'ha7, 8'hbb}; // CH=6 OP=1
cfg[2510] = { 1'b1, 8'hac, 8'h3b}; // CH=3 OP=3
cfg[2511] = { 1'b0, 8'h73, 8'hf9}; // CH=3 OP=0
cfg[2512] = { 1'b1, 8'he5, 8'h84}; // CH=4 OP=1
cfg[2513] = { 1'b0, 8'he2, 8'h43}; // CH=2 OP=0
cfg[2514] = { 1'b1, 8'h51, 8'h25}; // CH=4 OP=0
cfg[2515] = { 1'b1, 8'h67, 8'hef}; // CH=6 OP=1
cfg[2516] = { 1'b1, 8'hc0, 8'h12}; // CH=3 OP=0
cfg[2517] = { 1'b0, 8'hc9, 8'h1e}; // CH=1 OP=2
cfg[2518] = { 1'b1, 8'h84, 8'h10}; // CH=3 OP=1
cfg[2519] = { 1'b0, 8'hbf, 8'h8f}; // CH=3 OP=3
cfg[2520] = { 1'b0, 8'hb8, 8'hdd}; // CH=0 OP=2
cfg[2521] = { 1'b0, 8'h3c, 8'h5e}; // CH=0 OP=3
cfg[2522] = { 1'b1, 8'h7f, 8'hde}; // CH=6 OP=3
cfg[2523] = { 1'b0, 8'ha5, 8'he5}; // CH=1 OP=1
cfg[2524] = { 1'b1, 8'h94, 8'hc4}; // CH=3 OP=1
cfg[2525] = { 1'b1, 8'ha4, 8'h2c}; // CH=3 OP=1
cfg[2526] = { 1'b1, 8'hab, 8'h43}; // CH=6 OP=2
cfg[2527] = { 1'b0, 8'hc9, 8'h57}; // CH=1 OP=2
cfg[2528] = { 1'b1, 8'hd9, 8'h3a}; // CH=4 OP=2
cfg[2529] = { 1'b0, 8'h68, 8'hc4}; // CH=0 OP=2
cfg[2530] = { 1'b1, 8'h45, 8'hfb}; // CH=4 OP=1
cfg[2531] = { 1'b0, 8'ha3, 8'ha5}; // CH=3 OP=0
cfg[2532] = { 1'b0, 8'h81, 8'h34}; // CH=1 OP=0
cfg[2533] = { 1'b0, 8'h66, 8'ha6}; // CH=2 OP=1
cfg[2534] = { 1'b1, 8'h57, 8'h69}; // CH=6 OP=1
cfg[2535] = { 1'b1, 8'hfb, 8'h57}; // CH=6 OP=2
cfg[2536] = { 1'b0, 8'ha6, 8'h9a}; // CH=2 OP=1
cfg[2537] = { 1'b0, 8'h70, 8'hf1}; // CH=0 OP=0
cfg[2538] = { 1'b0, 8'h49, 8'h2c}; // CH=1 OP=2
cfg[2539] = { 1'b0, 8'hb2, 8'hf0}; // CH=2 OP=0
cfg[2540] = { 1'b1, 8'hf7, 8'heb}; // CH=6 OP=1
cfg[2541] = { 1'b1, 8'h9b, 8'h90}; // CH=6 OP=2
cfg[2542] = { 1'b0, 8'hc2, 8'hc5}; // CH=2 OP=0
cfg[2543] = { 1'b1, 8'h85, 8'h83}; // CH=4 OP=1
cfg[2544] = { 1'b1, 8'hdc, 8'hae}; // CH=3 OP=3
cfg[2545] = { 1'b0, 8'hd8, 8'h5}; // CH=0 OP=2
cfg[2546] = { 1'b0, 8'h7e, 8'h9f}; // CH=2 OP=3
cfg[2547] = { 1'b1, 8'hee, 8'h90}; // CH=5 OP=3
cfg[2548] = { 1'b1, 8'h38, 8'hbc}; // CH=3 OP=2
cfg[2549] = { 1'b1, 8'hea, 8'had}; // CH=5 OP=2
cfg[2550] = { 1'b0, 8'he1, 8'h98}; // CH=1 OP=0
cfg[2551] = { 1'b0, 8'h7c, 8'h29}; // CH=0 OP=3
cfg[2552] = { 1'b0, 8'h99, 8'hee}; // CH=1 OP=2
cfg[2553] = { 1'b0, 8'h5f, 8'h59}; // CH=3 OP=3
cfg[2554] = { 1'b0, 8'h3b, 8'hca}; // CH=3 OP=2
cfg[2555] = { 1'b0, 8'h4d, 8'hcf}; // CH=1 OP=3
cfg[2556] = { 1'b0, 8'hfe, 8'h92}; // CH=2 OP=3
cfg[2557] = { 1'b0, 8'hbb, 8'hdf}; // CH=3 OP=2
cfg[2558] = { 1'b0, 8'h68, 8'haa}; // CH=0 OP=2
cfg[2559] = { 1'b0, 8'h84, 8'h18}; // CH=0 OP=1
cfg[2560] = { 1'b0, 8'ha4, 8'h29}; // CH=0 OP=1
cfg[2561] = { 1'b1, 8'h7e, 8'h99}; // CH=5 OP=3
cfg[2562] = { 1'b1, 8'hdd, 8'hb5}; // CH=4 OP=3
cfg[2563] = { 1'b1, 8'hd6, 8'h7f}; // CH=5 OP=1
cfg[2564] = { 1'b0, 8'hbc, 8'h2c}; // CH=0 OP=3
cfg[2565] = { 1'b0, 8'hbb, 8'h31}; // CH=3 OP=2
cfg[2566] = { 1'b1, 8'h76, 8'h10}; // CH=5 OP=1
cfg[2567] = { 1'b1, 8'hde, 8'hba}; // CH=5 OP=3
cfg[2568] = { 1'b0, 8'hde, 8'hd2}; // CH=2 OP=3
cfg[2569] = { 1'b0, 8'hb8, 8'h5f}; // CH=0 OP=2
cfg[2570] = { 1'b0, 8'h6d, 8'h90}; // CH=1 OP=3
cfg[2571] = { 1'b1, 8'hed, 8'h30}; // CH=4 OP=3
cfg[2572] = { 1'b0, 8'h3b, 8'h6}; // CH=3 OP=2
cfg[2573] = { 1'b1, 8'hf8, 8'h29}; // CH=3 OP=2
cfg[2574] = { 1'b1, 8'hb3, 8'h5a}; // CH=6 OP=0
cfg[2575] = { 1'b0, 8'h9a, 8'h6a}; // CH=2 OP=2
cfg[2576] = { 1'b0, 8'h34, 8'h7}; // CH=0 OP=1
cfg[2577] = { 1'b0, 8'h52, 8'he5}; // CH=2 OP=0
cfg[2578] = { 1'b1, 8'h70, 8'hed}; // CH=3 OP=0
cfg[2579] = { 1'b1, 8'hdb, 8'hd}; // CH=6 OP=2
cfg[2580] = { 1'b1, 8'h3a, 8'h96}; // CH=5 OP=2
cfg[2581] = { 1'b1, 8'hb3, 8'h83}; // CH=6 OP=0
cfg[2582] = { 1'b1, 8'h58, 8'hbe}; // CH=3 OP=2
cfg[2583] = { 1'b0, 8'hbb, 8'hb6}; // CH=3 OP=2
cfg[2584] = { 1'b0, 8'h5e, 8'h69}; // CH=2 OP=3
cfg[2585] = { 1'b0, 8'hf8, 8'h92}; // CH=0 OP=2
cfg[2586] = { 1'b0, 8'hdb, 8'h99}; // CH=3 OP=2
cfg[2587] = { 1'b1, 8'h30, 8'h7e}; // CH=3 OP=0
cfg[2588] = { 1'b0, 8'h89, 8'hee}; // CH=1 OP=2
cfg[2589] = { 1'b1, 8'h64, 8'h17}; // CH=3 OP=1
cfg[2590] = { 1'b1, 8'h9f, 8'had}; // CH=6 OP=3
cfg[2591] = { 1'b0, 8'h52, 8'h30}; // CH=2 OP=0
cfg[2592] = { 1'b0, 8'haa, 8'hee}; // CH=2 OP=2
cfg[2593] = { 1'b0, 8'h65, 8'ha5}; // CH=1 OP=1
cfg[2594] = { 1'b1, 8'hc3, 8'he}; // CH=6 OP=0
cfg[2595] = { 1'b1, 8'hbb, 8'ha1}; // CH=6 OP=2
cfg[2596] = { 1'b0, 8'he7, 8'h3a}; // CH=3 OP=1
cfg[2597] = { 1'b1, 8'h65, 8'hb9}; // CH=4 OP=1
cfg[2598] = { 1'b1, 8'h54, 8'h26}; // CH=3 OP=1
cfg[2599] = { 1'b1, 8'h6b, 8'h9f}; // CH=6 OP=2
cfg[2600] = { 1'b1, 8'h48, 8'hb6}; // CH=3 OP=2
cfg[2601] = { 1'b1, 8'h9a, 8'h48}; // CH=5 OP=2
cfg[2602] = { 1'b1, 8'h44, 8'h36}; // CH=3 OP=1
cfg[2603] = { 1'b1, 8'haa, 8'hdb}; // CH=5 OP=2
cfg[2604] = { 1'b0, 8'h6d, 8'hea}; // CH=1 OP=3
cfg[2605] = { 1'b0, 8'h8e, 8'h8b}; // CH=2 OP=3
cfg[2606] = { 1'b1, 8'h7f, 8'h10}; // CH=6 OP=3
cfg[2607] = { 1'b0, 8'ha5, 8'hd4}; // CH=1 OP=1
cfg[2608] = { 1'b0, 8'h44, 8'h19}; // CH=0 OP=1
cfg[2609] = { 1'b1, 8'hfb, 8'hc3}; // CH=6 OP=2
cfg[2610] = { 1'b1, 8'h96, 8'hb}; // CH=5 OP=1
cfg[2611] = { 1'b1, 8'he9, 8'ha6}; // CH=4 OP=2
cfg[2612] = { 1'b1, 8'hf0, 8'hea}; // CH=3 OP=0
cfg[2613] = { 1'b1, 8'h91, 8'h94}; // CH=4 OP=0
cfg[2614] = { 1'b0, 8'h6f, 8'he1}; // CH=3 OP=3
cfg[2615] = { 1'b1, 8'h88, 8'h3b}; // CH=3 OP=2
cfg[2616] = { 1'b0, 8'h5c, 8'hb1}; // CH=0 OP=3
cfg[2617] = { 1'b1, 8'h76, 8'h7b}; // CH=5 OP=1
cfg[2618] = { 1'b0, 8'h39, 8'hb0}; // CH=1 OP=2
cfg[2619] = { 1'b1, 8'h44, 8'hfd}; // CH=3 OP=1
cfg[2620] = { 1'b1, 8'hea, 8'h92}; // CH=5 OP=2
cfg[2621] = { 1'b0, 8'hd5, 8'h5e}; // CH=1 OP=1
cfg[2622] = { 1'b0, 8'h69, 8'h5}; // CH=1 OP=2
cfg[2623] = { 1'b1, 8'h6b, 8'h96}; // CH=6 OP=2
cfg[2624] = { 1'b0, 8'h96, 8'hb2}; // CH=2 OP=1
cfg[2625] = { 1'b1, 8'hd2, 8'h93}; // CH=5 OP=0
cfg[2626] = { 1'b1, 8'h83, 8'hf4}; // CH=6 OP=0
cfg[2627] = { 1'b0, 8'hff, 8'hf9}; // CH=3 OP=3
cfg[2628] = { 1'b0, 8'haf, 8'h43}; // CH=3 OP=3
cfg[2629] = { 1'b1, 8'had, 8'h88}; // CH=4 OP=3
cfg[2630] = { 1'b1, 8'h3f, 8'h63}; // CH=6 OP=3
cfg[2631] = { 1'b0, 8'h9d, 8'h27}; // CH=1 OP=3
cfg[2632] = { 1'b1, 8'ha2, 8'hdc}; // CH=5 OP=0
cfg[2633] = { 1'b0, 8'h38, 8'h93}; // CH=0 OP=2
cfg[2634] = { 1'b0, 8'hea, 8'h2c}; // CH=2 OP=2
cfg[2635] = { 1'b0, 8'h7e, 8'h33}; // CH=2 OP=3
cfg[2636] = { 1'b0, 8'h72, 8'hc3}; // CH=2 OP=0
cfg[2637] = { 1'b0, 8'h6b, 8'haf}; // CH=3 OP=2
cfg[2638] = { 1'b1, 8'haf, 8'h11}; // CH=6 OP=3
cfg[2639] = { 1'b0, 8'h37, 8'hac}; // CH=3 OP=1
cfg[2640] = { 1'b1, 8'h9b, 8'h8b}; // CH=6 OP=2
cfg[2641] = { 1'b1, 8'hc2, 8'h55}; // CH=5 OP=0
cfg[2642] = { 1'b0, 8'h9e, 8'hf4}; // CH=2 OP=3
cfg[2643] = { 1'b1, 8'h32, 8'hfd}; // CH=5 OP=0
cfg[2644] = { 1'b1, 8'h5e, 8'h71}; // CH=5 OP=3
cfg[2645] = { 1'b0, 8'h91, 8'h7b}; // CH=1 OP=0
cfg[2646] = { 1'b0, 8'h54, 8'h58}; // CH=0 OP=1
cfg[2647] = { 1'b0, 8'hb9, 8'hb8}; // CH=1 OP=2
cfg[2648] = { 1'b1, 8'h68, 8'h14}; // CH=3 OP=2
cfg[2649] = { 1'b1, 8'ha0, 8'hc0}; // CH=3 OP=0
cfg[2650] = { 1'b1, 8'h3b, 8'h4c}; // CH=6 OP=2
cfg[2651] = { 1'b0, 8'hfd, 8'ha1}; // CH=1 OP=3
cfg[2652] = { 1'b0, 8'h9c, 8'h96}; // CH=0 OP=3
cfg[2653] = { 1'b1, 8'hce, 8'h93}; // CH=5 OP=3
cfg[2654] = { 1'b1, 8'h81, 8'h4}; // CH=4 OP=0
cfg[2655] = { 1'b1, 8'h5d, 8'hbd}; // CH=4 OP=3
cfg[2656] = { 1'b1, 8'hab, 8'h12}; // CH=6 OP=2
cfg[2657] = { 1'b1, 8'h64, 8'h15}; // CH=3 OP=1
cfg[2658] = { 1'b0, 8'hcd, 8'h2a}; // CH=1 OP=3
cfg[2659] = { 1'b0, 8'h6d, 8'hea}; // CH=1 OP=3
cfg[2660] = { 1'b1, 8'ha8, 8'h36}; // CH=3 OP=2
cfg[2661] = { 1'b1, 8'ha5, 8'hd8}; // CH=4 OP=1
cfg[2662] = { 1'b1, 8'h41, 8'h6e}; // CH=4 OP=0
cfg[2663] = { 1'b1, 8'hd0, 8'h1}; // CH=3 OP=0
cfg[2664] = { 1'b1, 8'h51, 8'h3b}; // CH=4 OP=0
cfg[2665] = { 1'b0, 8'hae, 8'hf9}; // CH=2 OP=3
cfg[2666] = { 1'b0, 8'h59, 8'hb}; // CH=1 OP=2
cfg[2667] = { 1'b1, 8'hbd, 8'h20}; // CH=4 OP=3
cfg[2668] = { 1'b0, 8'h8a, 8'h4a}; // CH=2 OP=2
cfg[2669] = { 1'b0, 8'hf7, 8'h35}; // CH=3 OP=1
cfg[2670] = { 1'b1, 8'h9f, 8'h6b}; // CH=6 OP=3
cfg[2671] = { 1'b0, 8'h45, 8'h43}; // CH=1 OP=1
cfg[2672] = { 1'b1, 8'h86, 8'hb1}; // CH=5 OP=1
cfg[2673] = { 1'b0, 8'h96, 8'hb2}; // CH=2 OP=1
cfg[2674] = { 1'b0, 8'hd1, 8'hb7}; // CH=1 OP=0
cfg[2675] = { 1'b1, 8'hca, 8'h3c}; // CH=5 OP=2
cfg[2676] = { 1'b1, 8'hd5, 8'h98}; // CH=4 OP=1
cfg[2677] = { 1'b0, 8'hf6, 8'h83}; // CH=2 OP=1
cfg[2678] = { 1'b0, 8'h40, 8'h15}; // CH=0 OP=0
cfg[2679] = { 1'b0, 8'h75, 8'h73}; // CH=1 OP=1
cfg[2680] = { 1'b0, 8'he1, 8'h7e}; // CH=1 OP=0
cfg[2681] = { 1'b1, 8'h8a, 8'h12}; // CH=5 OP=2
cfg[2682] = { 1'b0, 8'he2, 8'hd6}; // CH=2 OP=0
cfg[2683] = { 1'b0, 8'hf1, 8'ha7}; // CH=1 OP=0
cfg[2684] = { 1'b0, 8'h50, 8'h78}; // CH=0 OP=0
cfg[2685] = { 1'b0, 8'h5e, 8'h43}; // CH=2 OP=3
cfg[2686] = { 1'b0, 8'hc4, 8'h18}; // CH=0 OP=1
cfg[2687] = { 1'b1, 8'he8, 8'he}; // CH=3 OP=2
cfg[2688] = { 1'b1, 8'h97, 8'h4f}; // CH=6 OP=1
cfg[2689] = { 1'b0, 8'h3d, 8'hc4}; // CH=1 OP=3
cfg[2690] = { 1'b1, 8'h82, 8'ha5}; // CH=5 OP=0
cfg[2691] = { 1'b1, 8'h55, 8'hca}; // CH=4 OP=1
cfg[2692] = { 1'b0, 8'h38, 8'h1e}; // CH=0 OP=2
cfg[2693] = { 1'b0, 8'h68, 8'hc5}; // CH=0 OP=2
cfg[2694] = { 1'b1, 8'he4, 8'h79}; // CH=3 OP=1
cfg[2695] = { 1'b0, 8'hf8, 8'hd7}; // CH=0 OP=2
cfg[2696] = { 1'b1, 8'h90, 8'h9c}; // CH=3 OP=0
cfg[2697] = { 1'b1, 8'h3d, 8'h84}; // CH=4 OP=3
cfg[2698] = { 1'b0, 8'h5d, 8'h1b}; // CH=1 OP=3
cfg[2699] = { 1'b1, 8'hfc, 8'h58}; // CH=3 OP=3
cfg[2700] = { 1'b0, 8'hae, 8'hdb}; // CH=2 OP=3
cfg[2701] = { 1'b0, 8'hca, 8'he8}; // CH=2 OP=2
cfg[2702] = { 1'b0, 8'hf3, 8'h3b}; // CH=3 OP=0
cfg[2703] = { 1'b1, 8'h5b, 8'h64}; // CH=6 OP=2
cfg[2704] = { 1'b0, 8'h40, 8'hde}; // CH=0 OP=0
cfg[2705] = { 1'b1, 8'h38, 8'hb5}; // CH=3 OP=2
cfg[2706] = { 1'b0, 8'hc8, 8'h51}; // CH=0 OP=2
cfg[2707] = { 1'b1, 8'hc0, 8'hd6}; // CH=3 OP=0
cfg[2708] = { 1'b1, 8'h7b, 8'h63}; // CH=6 OP=2
cfg[2709] = { 1'b0, 8'hdb, 8'h5f}; // CH=3 OP=2
cfg[2710] = { 1'b1, 8'hd0, 8'hd}; // CH=3 OP=0
cfg[2711] = { 1'b1, 8'hc3, 8'h4c}; // CH=6 OP=0
cfg[2712] = { 1'b0, 8'he6, 8'hb1}; // CH=2 OP=1
cfg[2713] = { 1'b1, 8'h6f, 8'h5f}; // CH=6 OP=3
cfg[2714] = { 1'b0, 8'h91, 8'h97}; // CH=1 OP=0
cfg[2715] = { 1'b0, 8'h5b, 8'h60}; // CH=3 OP=2
cfg[2716] = { 1'b0, 8'h5d, 8'h65}; // CH=1 OP=3
cfg[2717] = { 1'b0, 8'ha7, 8'h96}; // CH=3 OP=1
cfg[2718] = { 1'b0, 8'hcc, 8'h71}; // CH=0 OP=3
cfg[2719] = { 1'b1, 8'hd9, 8'h77}; // CH=4 OP=2
cfg[2720] = { 1'b0, 8'hec, 8'h48}; // CH=0 OP=3
cfg[2721] = { 1'b1, 8'hca, 8'hb}; // CH=5 OP=2
cfg[2722] = { 1'b0, 8'hb1, 8'h2a}; // CH=1 OP=0
cfg[2723] = { 1'b1, 8'hb2, 8'h89}; // CH=5 OP=0
cfg[2724] = { 1'b1, 8'he6, 8'h81}; // CH=5 OP=1
cfg[2725] = { 1'b0, 8'haf, 8'h77}; // CH=3 OP=3
cfg[2726] = { 1'b0, 8'hd7, 8'h1e}; // CH=3 OP=1
cfg[2727] = { 1'b1, 8'ha7, 8'heb}; // CH=6 OP=1
cfg[2728] = { 1'b0, 8'hef, 8'h53}; // CH=3 OP=3
cfg[2729] = { 1'b1, 8'hfa, 8'he6}; // CH=5 OP=2
cfg[2730] = { 1'b1, 8'hfd, 8'h2a}; // CH=4 OP=3
cfg[2731] = { 1'b0, 8'hcf, 8'h4d}; // CH=3 OP=3
cfg[2732] = { 1'b1, 8'h50, 8'hc2}; // CH=3 OP=0
cfg[2733] = { 1'b0, 8'h37, 8'hdb}; // CH=3 OP=1
cfg[2734] = { 1'b0, 8'he6, 8'h52}; // CH=2 OP=1
cfg[2735] = { 1'b0, 8'hbd, 8'h71}; // CH=1 OP=3
cfg[2736] = { 1'b1, 8'hc9, 8'h5c}; // CH=4 OP=2
cfg[2737] = { 1'b0, 8'hb7, 8'h20}; // CH=3 OP=1
cfg[2738] = { 1'b1, 8'hb2, 8'h2}; // CH=5 OP=0
cfg[2739] = { 1'b1, 8'hd7, 8'h2c}; // CH=6 OP=1
cfg[2740] = { 1'b1, 8'h85, 8'h29}; // CH=4 OP=1
cfg[2741] = { 1'b0, 8'h55, 8'h3e}; // CH=1 OP=1
cfg[2742] = { 1'b1, 8'ha5, 8'h0}; // CH=4 OP=1
cfg[2743] = { 1'b1, 8'hdc, 8'hdb}; // CH=3 OP=3
cfg[2744] = { 1'b1, 8'hc2, 8'h2e}; // CH=5 OP=0
cfg[2745] = { 1'b1, 8'h7f, 8'h9f}; // CH=6 OP=3
cfg[2746] = { 1'b1, 8'h49, 8'hfb}; // CH=4 OP=2
cfg[2747] = { 1'b1, 8'h65, 8'h1b}; // CH=4 OP=1
cfg[2748] = { 1'b1, 8'h68, 8'hed}; // CH=3 OP=2
cfg[2749] = { 1'b1, 8'h94, 8'h3a}; // CH=3 OP=1
cfg[2750] = { 1'b0, 8'hbe, 8'hb3}; // CH=2 OP=3
cfg[2751] = { 1'b1, 8'hfc, 8'h7a}; // CH=3 OP=3
cfg[2752] = { 1'b0, 8'hfc, 8'h3f}; // CH=0 OP=3
cfg[2753] = { 1'b0, 8'hd7, 8'h11}; // CH=3 OP=1
cfg[2754] = { 1'b0, 8'h41, 8'h16}; // CH=1 OP=0
cfg[2755] = { 1'b0, 8'hc0, 8'ha4}; // CH=0 OP=0
cfg[2756] = { 1'b1, 8'hbb, 8'h9f}; // CH=6 OP=2
cfg[2757] = { 1'b1, 8'ha8, 8'ha1}; // CH=3 OP=2
cfg[2758] = { 1'b1, 8'he2, 8'hec}; // CH=5 OP=0
cfg[2759] = { 1'b1, 8'h95, 8'he}; // CH=4 OP=1
cfg[2760] = { 1'b1, 8'hb2, 8'hb6}; // CH=5 OP=0
cfg[2761] = { 1'b1, 8'h54, 8'h21}; // CH=3 OP=1
cfg[2762] = { 1'b0, 8'hd3, 8'hf9}; // CH=3 OP=0
cfg[2763] = { 1'b0, 8'h84, 8'hfe}; // CH=0 OP=1
cfg[2764] = { 1'b1, 8'hab, 8'hd4}; // CH=6 OP=2
cfg[2765] = { 1'b0, 8'hb4, 8'hde}; // CH=0 OP=1
cfg[2766] = { 1'b1, 8'h55, 8'h4d}; // CH=4 OP=1
cfg[2767] = { 1'b1, 8'h42, 8'h24}; // CH=5 OP=0
cfg[2768] = { 1'b1, 8'h50, 8'h8f}; // CH=3 OP=0
cfg[2769] = { 1'b1, 8'hde, 8'hb9}; // CH=5 OP=3
cfg[2770] = { 1'b1, 8'hdb, 8'h7b}; // CH=6 OP=2
cfg[2771] = { 1'b1, 8'h52, 8'he0}; // CH=5 OP=0
cfg[2772] = { 1'b1, 8'hd6, 8'hf4}; // CH=5 OP=1
cfg[2773] = { 1'b0, 8'h82, 8'hc9}; // CH=2 OP=0
cfg[2774] = { 1'b1, 8'h36, 8'ha7}; // CH=5 OP=1
cfg[2775] = { 1'b0, 8'h8b, 8'hf4}; // CH=3 OP=2
cfg[2776] = { 1'b0, 8'hcd, 8'h18}; // CH=1 OP=3
cfg[2777] = { 1'b1, 8'h60, 8'ha7}; // CH=3 OP=0
cfg[2778] = { 1'b0, 8'h3f, 8'h51}; // CH=3 OP=3
cfg[2779] = { 1'b1, 8'h3f, 8'hcc}; // CH=6 OP=3
cfg[2780] = { 1'b1, 8'h38, 8'ha8}; // CH=3 OP=2
cfg[2781] = { 1'b1, 8'hc0, 8'hfa}; // CH=3 OP=0
cfg[2782] = { 1'b0, 8'h89, 8'hca}; // CH=1 OP=2
cfg[2783] = { 1'b0, 8'h30, 8'ha7}; // CH=0 OP=0
cfg[2784] = { 1'b0, 8'h3c, 8'h81}; // CH=0 OP=3
cfg[2785] = { 1'b1, 8'he3, 8'h9}; // CH=6 OP=0
cfg[2786] = { 1'b1, 8'h44, 8'h2d}; // CH=3 OP=1
cfg[2787] = { 1'b0, 8'h83, 8'h7e}; // CH=3 OP=0
cfg[2788] = { 1'b1, 8'hc2, 8'h4b}; // CH=5 OP=0
cfg[2789] = { 1'b0, 8'hfa, 8'hf3}; // CH=2 OP=2
cfg[2790] = { 1'b0, 8'h78, 8'hed}; // CH=0 OP=2
cfg[2791] = { 1'b1, 8'h9a, 8'hf3}; // CH=5 OP=2
cfg[2792] = { 1'b1, 8'h55, 8'h98}; // CH=4 OP=1
cfg[2793] = { 1'b0, 8'h91, 8'h1d}; // CH=1 OP=0
cfg[2794] = { 1'b0, 8'h74, 8'h26}; // CH=0 OP=1
cfg[2795] = { 1'b1, 8'hb8, 8'h54}; // CH=3 OP=2
cfg[2796] = { 1'b1, 8'h3b, 8'hd2}; // CH=6 OP=2
cfg[2797] = { 1'b1, 8'hfd, 8'h1d}; // CH=4 OP=3
cfg[2798] = { 1'b1, 8'hf7, 8'h10}; // CH=6 OP=1
cfg[2799] = { 1'b1, 8'hcf, 8'hfd}; // CH=6 OP=3
cfg[2800] = { 1'b1, 8'hd0, 8'h14}; // CH=3 OP=0
cfg[2801] = { 1'b1, 8'h63, 8'haf}; // CH=6 OP=0
cfg[2802] = { 1'b1, 8'he8, 8'h56}; // CH=3 OP=2
cfg[2803] = { 1'b1, 8'h5c, 8'h9e}; // CH=3 OP=3
cfg[2804] = { 1'b1, 8'hdd, 8'h63}; // CH=4 OP=3
cfg[2805] = { 1'b1, 8'h90, 8'h50}; // CH=3 OP=0
cfg[2806] = { 1'b1, 8'h63, 8'h4d}; // CH=6 OP=0
cfg[2807] = { 1'b1, 8'h61, 8'h87}; // CH=4 OP=0
cfg[2808] = { 1'b0, 8'h7a, 8'h56}; // CH=2 OP=2
cfg[2809] = { 1'b1, 8'h4a, 8'he7}; // CH=5 OP=2
cfg[2810] = { 1'b0, 8'h5a, 8'h7f}; // CH=2 OP=2
cfg[2811] = { 1'b1, 8'hf8, 8'h66}; // CH=3 OP=2
cfg[2812] = { 1'b0, 8'h4f, 8'hc2}; // CH=3 OP=3
cfg[2813] = { 1'b1, 8'h84, 8'h1}; // CH=3 OP=1
cfg[2814] = { 1'b1, 8'hd7, 8'h91}; // CH=6 OP=1
cfg[2815] = { 1'b0, 8'h3b, 8'hc0}; // CH=3 OP=2
cfg[2816] = { 1'b1, 8'h9c, 8'h47}; // CH=3 OP=3
cfg[2817] = { 1'b1, 8'hb8, 8'h9e}; // CH=3 OP=2
cfg[2818] = { 1'b0, 8'h9f, 8'hc5}; // CH=3 OP=3
cfg[2819] = { 1'b1, 8'he9, 8'hed}; // CH=4 OP=2
cfg[2820] = { 1'b0, 8'h44, 8'h6c}; // CH=0 OP=1
cfg[2821] = { 1'b1, 8'h3c, 8'hd3}; // CH=3 OP=3
cfg[2822] = { 1'b1, 8'h60, 8'h95}; // CH=3 OP=0
cfg[2823] = { 1'b0, 8'h61, 8'h6c}; // CH=1 OP=0
cfg[2824] = { 1'b0, 8'hf2, 8'h93}; // CH=2 OP=0
cfg[2825] = { 1'b0, 8'hb3, 8'h8}; // CH=3 OP=0
cfg[2826] = { 1'b1, 8'hfa, 8'hc1}; // CH=5 OP=2
cfg[2827] = { 1'b1, 8'h98, 8'he1}; // CH=3 OP=2
cfg[2828] = { 1'b1, 8'h5d, 8'h7b}; // CH=4 OP=3
cfg[2829] = { 1'b0, 8'h4b, 8'h3e}; // CH=3 OP=2
cfg[2830] = { 1'b1, 8'hb7, 8'hf6}; // CH=6 OP=1
cfg[2831] = { 1'b1, 8'h8a, 8'h8b}; // CH=5 OP=2
cfg[2832] = { 1'b0, 8'hdc, 8'hc}; // CH=0 OP=3
cfg[2833] = { 1'b0, 8'h31, 8'h86}; // CH=1 OP=0
cfg[2834] = { 1'b0, 8'h5d, 8'h78}; // CH=1 OP=3
cfg[2835] = { 1'b0, 8'hc4, 8'h2b}; // CH=0 OP=1
cfg[2836] = { 1'b1, 8'hc7, 8'h26}; // CH=6 OP=1
cfg[2837] = { 1'b0, 8'h82, 8'hbe}; // CH=2 OP=0
cfg[2838] = { 1'b1, 8'hdc, 8'h1c}; // CH=3 OP=3
cfg[2839] = { 1'b0, 8'h7a, 8'h67}; // CH=2 OP=2
cfg[2840] = { 1'b0, 8'ha9, 8'ha7}; // CH=1 OP=2
cfg[2841] = { 1'b1, 8'hc9, 8'h12}; // CH=4 OP=2
cfg[2842] = { 1'b1, 8'h55, 8'hef}; // CH=4 OP=1
cfg[2843] = { 1'b1, 8'h75, 8'h20}; // CH=4 OP=1
cfg[2844] = { 1'b0, 8'h9d, 8'h7d}; // CH=1 OP=3
cfg[2845] = { 1'b1, 8'h87, 8'h41}; // CH=6 OP=1
cfg[2846] = { 1'b1, 8'h51, 8'h8}; // CH=4 OP=0
cfg[2847] = { 1'b0, 8'h97, 8'h8a}; // CH=3 OP=1
cfg[2848] = { 1'b0, 8'h85, 8'h66}; // CH=1 OP=1
cfg[2849] = { 1'b1, 8'h9b, 8'h3f}; // CH=6 OP=2
cfg[2850] = { 1'b0, 8'hae, 8'h97}; // CH=2 OP=3
cfg[2851] = { 1'b1, 8'h9d, 8'h27}; // CH=4 OP=3
cfg[2852] = { 1'b1, 8'hbd, 8'h3c}; // CH=4 OP=3
cfg[2853] = { 1'b0, 8'h3a, 8'hca}; // CH=2 OP=2
cfg[2854] = { 1'b0, 8'h7b, 8'h84}; // CH=3 OP=2
cfg[2855] = { 1'b1, 8'h83, 8'h63}; // CH=6 OP=0
cfg[2856] = { 1'b0, 8'h89, 8'h1}; // CH=1 OP=2
cfg[2857] = { 1'b1, 8'ha4, 8'h73}; // CH=3 OP=1
cfg[2858] = { 1'b0, 8'h3a, 8'hf8}; // CH=2 OP=2
cfg[2859] = { 1'b0, 8'hd5, 8'h25}; // CH=1 OP=1
cfg[2860] = { 1'b0, 8'h83, 8'hbc}; // CH=3 OP=0
cfg[2861] = { 1'b0, 8'hbd, 8'he3}; // CH=1 OP=3
cfg[2862] = { 1'b0, 8'h39, 8'hdd}; // CH=1 OP=2
cfg[2863] = { 1'b0, 8'h53, 8'h17}; // CH=3 OP=0
cfg[2864] = { 1'b0, 8'hf4, 8'h92}; // CH=0 OP=1
cfg[2865] = { 1'b0, 8'he7, 8'h15}; // CH=3 OP=1
cfg[2866] = { 1'b1, 8'h70, 8'h22}; // CH=3 OP=0
cfg[2867] = { 1'b1, 8'h6b, 8'h95}; // CH=6 OP=2
cfg[2868] = { 1'b0, 8'h87, 8'h4f}; // CH=3 OP=1
cfg[2869] = { 1'b1, 8'h8c, 8'h24}; // CH=3 OP=3
cfg[2870] = { 1'b1, 8'h42, 8'ha8}; // CH=5 OP=0
cfg[2871] = { 1'b1, 8'hff, 8'hc8}; // CH=6 OP=3
cfg[2872] = { 1'b1, 8'h38, 8'ha6}; // CH=3 OP=2
cfg[2873] = { 1'b1, 8'h8c, 8'hbd}; // CH=3 OP=3
cfg[2874] = { 1'b0, 8'h80, 8'h50}; // CH=0 OP=0
cfg[2875] = { 1'b0, 8'h67, 8'h65}; // CH=3 OP=1
cfg[2876] = { 1'b1, 8'hd8, 8'h88}; // CH=3 OP=2
cfg[2877] = { 1'b0, 8'hed, 8'h1d}; // CH=1 OP=3
cfg[2878] = { 1'b0, 8'h3c, 8'hab}; // CH=0 OP=3
cfg[2879] = { 1'b1, 8'h60, 8'h5e}; // CH=3 OP=0
cfg[2880] = { 1'b1, 8'hc1, 8'hce}; // CH=4 OP=0
cfg[2881] = { 1'b1, 8'hc0, 8'hd1}; // CH=3 OP=0
cfg[2882] = { 1'b0, 8'hf9, 8'h77}; // CH=1 OP=2
cfg[2883] = { 1'b1, 8'h85, 8'h34}; // CH=4 OP=1
cfg[2884] = { 1'b1, 8'h5b, 8'h84}; // CH=6 OP=2
cfg[2885] = { 1'b0, 8'hcd, 8'h6d}; // CH=1 OP=3
cfg[2886] = { 1'b0, 8'hcd, 8'h45}; // CH=1 OP=3
cfg[2887] = { 1'b1, 8'h39, 8'h32}; // CH=4 OP=2
cfg[2888] = { 1'b1, 8'h99, 8'h6e}; // CH=4 OP=2
cfg[2889] = { 1'b0, 8'h67, 8'hac}; // CH=3 OP=1
cfg[2890] = { 1'b1, 8'h88, 8'h6e}; // CH=3 OP=2
cfg[2891] = { 1'b0, 8'h53, 8'h2e}; // CH=3 OP=0
cfg[2892] = { 1'b0, 8'hd8, 8'hcb}; // CH=0 OP=2
cfg[2893] = { 1'b0, 8'hc2, 8'h27}; // CH=2 OP=0
cfg[2894] = { 1'b1, 8'h34, 8'hf4}; // CH=3 OP=1
cfg[2895] = { 1'b0, 8'hc3, 8'hc1}; // CH=3 OP=0
cfg[2896] = { 1'b0, 8'hfe, 8'hfb}; // CH=2 OP=3
cfg[2897] = { 1'b0, 8'h98, 8'h28}; // CH=0 OP=2
cfg[2898] = { 1'b0, 8'hff, 8'hd4}; // CH=3 OP=3
cfg[2899] = { 1'b1, 8'h88, 8'h42}; // CH=3 OP=2
cfg[2900] = { 1'b1, 8'ha4, 8'h71}; // CH=3 OP=1
cfg[2901] = { 1'b0, 8'hb2, 8'h98}; // CH=2 OP=0
cfg[2902] = { 1'b0, 8'h7e, 8'h45}; // CH=2 OP=3
cfg[2903] = { 1'b0, 8'ha5, 8'hf7}; // CH=1 OP=1
cfg[2904] = { 1'b0, 8'h99, 8'h16}; // CH=1 OP=2
cfg[2905] = { 1'b0, 8'h5a, 8'h7a}; // CH=2 OP=2
cfg[2906] = { 1'b1, 8'h55, 8'h10}; // CH=4 OP=1
cfg[2907] = { 1'b0, 8'h7d, 8'h14}; // CH=1 OP=3
cfg[2908] = { 1'b0, 8'h52, 8'he6}; // CH=2 OP=0
cfg[2909] = { 1'b1, 8'h94, 8'h90}; // CH=3 OP=1
cfg[2910] = { 1'b1, 8'h52, 8'he1}; // CH=5 OP=0
cfg[2911] = { 1'b0, 8'he3, 8'hca}; // CH=3 OP=0
cfg[2912] = { 1'b0, 8'hda, 8'hb2}; // CH=2 OP=2
cfg[2913] = { 1'b1, 8'hf0, 8'h10}; // CH=3 OP=0
cfg[2914] = { 1'b0, 8'h6a, 8'ha2}; // CH=2 OP=2
cfg[2915] = { 1'b1, 8'h7a, 8'hf7}; // CH=5 OP=2
cfg[2916] = { 1'b0, 8'h8e, 8'h4b}; // CH=2 OP=3
cfg[2917] = { 1'b0, 8'h74, 8'h37}; // CH=0 OP=1
cfg[2918] = { 1'b0, 8'h9a, 8'h23}; // CH=2 OP=2
cfg[2919] = { 1'b0, 8'ha0, 8'he6}; // CH=0 OP=0
cfg[2920] = { 1'b0, 8'h3e, 8'h38}; // CH=2 OP=3
cfg[2921] = { 1'b1, 8'hc1, 8'h4e}; // CH=4 OP=0
cfg[2922] = { 1'b0, 8'haf, 8'hfb}; // CH=3 OP=3
cfg[2923] = { 1'b0, 8'h35, 8'heb}; // CH=1 OP=1
cfg[2924] = { 1'b0, 8'ha9, 8'h55}; // CH=1 OP=2
cfg[2925] = { 1'b1, 8'hf5, 8'h4d}; // CH=4 OP=1
cfg[2926] = { 1'b1, 8'hd1, 8'h1}; // CH=4 OP=0
cfg[2927] = { 1'b1, 8'hd6, 8'h4f}; // CH=5 OP=1
cfg[2928] = { 1'b1, 8'hbc, 8'he6}; // CH=3 OP=3
cfg[2929] = { 1'b1, 8'hf4, 8'h94}; // CH=3 OP=1
cfg[2930] = { 1'b1, 8'h42, 8'hd}; // CH=5 OP=0
cfg[2931] = { 1'b0, 8'h42, 8'hcf}; // CH=2 OP=0
cfg[2932] = { 1'b1, 8'h52, 8'h7e}; // CH=5 OP=0
cfg[2933] = { 1'b0, 8'hdb, 8'hb3}; // CH=3 OP=2
cfg[2934] = { 1'b0, 8'haa, 8'had}; // CH=2 OP=2
cfg[2935] = { 1'b1, 8'hcf, 8'ha2}; // CH=6 OP=3
cfg[2936] = { 1'b1, 8'haf, 8'h1f}; // CH=6 OP=3
cfg[2937] = { 1'b0, 8'h6b, 8'h4}; // CH=3 OP=2
cfg[2938] = { 1'b0, 8'h5f, 8'h99}; // CH=3 OP=3
cfg[2939] = { 1'b1, 8'ha1, 8'ha6}; // CH=4 OP=0
cfg[2940] = { 1'b0, 8'he3, 8'h75}; // CH=3 OP=0
cfg[2941] = { 1'b1, 8'h35, 8'hf3}; // CH=4 OP=1
cfg[2942] = { 1'b0, 8'h39, 8'ha7}; // CH=1 OP=2
cfg[2943] = { 1'b1, 8'he6, 8'h71}; // CH=5 OP=1
cfg[2944] = { 1'b0, 8'h89, 8'h88}; // CH=1 OP=2
cfg[2945] = { 1'b1, 8'h58, 8'ha0}; // CH=3 OP=2
cfg[2946] = { 1'b0, 8'h76, 8'hbf}; // CH=2 OP=1
cfg[2947] = { 1'b1, 8'h7b, 8'h7f}; // CH=6 OP=2
cfg[2948] = { 1'b0, 8'hba, 8'h81}; // CH=2 OP=2
cfg[2949] = { 1'b0, 8'h30, 8'h25}; // CH=0 OP=0
cfg[2950] = { 1'b1, 8'hdc, 8'he2}; // CH=3 OP=3
cfg[2951] = { 1'b0, 8'h46, 8'hca}; // CH=2 OP=1
cfg[2952] = { 1'b1, 8'hc3, 8'hfc}; // CH=6 OP=0
cfg[2953] = { 1'b1, 8'h63, 8'he1}; // CH=6 OP=0
cfg[2954] = { 1'b1, 8'h53, 8'h8c}; // CH=6 OP=0
cfg[2955] = { 1'b1, 8'hce, 8'ha2}; // CH=5 OP=3
cfg[2956] = { 1'b0, 8'he2, 8'h23}; // CH=2 OP=0
cfg[2957] = { 1'b1, 8'h9d, 8'h26}; // CH=4 OP=3
cfg[2958] = { 1'b0, 8'hcd, 8'h4b}; // CH=1 OP=3
cfg[2959] = { 1'b1, 8'hf0, 8'h2e}; // CH=3 OP=0
cfg[2960] = { 1'b0, 8'hbb, 8'h54}; // CH=3 OP=2
cfg[2961] = { 1'b1, 8'hf6, 8'h9a}; // CH=5 OP=1
cfg[2962] = { 1'b1, 8'hba, 8'haa}; // CH=5 OP=2
cfg[2963] = { 1'b0, 8'h89, 8'h8c}; // CH=1 OP=2
cfg[2964] = { 1'b0, 8'hdd, 8'h40}; // CH=1 OP=3
cfg[2965] = { 1'b1, 8'hab, 8'he2}; // CH=6 OP=2
cfg[2966] = { 1'b1, 8'h8e, 8'h5}; // CH=5 OP=3
cfg[2967] = { 1'b1, 8'h77, 8'h2c}; // CH=6 OP=1
cfg[2968] = { 1'b0, 8'ha5, 8'h40}; // CH=1 OP=1
cfg[2969] = { 1'b0, 8'hfa, 8'h56}; // CH=2 OP=2
cfg[2970] = { 1'b1, 8'h94, 8'h82}; // CH=3 OP=1
cfg[2971] = { 1'b0, 8'h3f, 8'ha9}; // CH=3 OP=3
cfg[2972] = { 1'b0, 8'hcb, 8'h56}; // CH=3 OP=2
cfg[2973] = { 1'b1, 8'he3, 8'hdf}; // CH=6 OP=0
cfg[2974] = { 1'b1, 8'he0, 8'hbc}; // CH=3 OP=0
cfg[2975] = { 1'b1, 8'h88, 8'h68}; // CH=3 OP=2
cfg[2976] = { 1'b1, 8'hfd, 8'hf6}; // CH=4 OP=3
cfg[2977] = { 1'b1, 8'h3c, 8'h21}; // CH=3 OP=3
cfg[2978] = { 1'b1, 8'he2, 8'h44}; // CH=5 OP=0
cfg[2979] = { 1'b1, 8'hdc, 8'h9b}; // CH=3 OP=3
cfg[2980] = { 1'b1, 8'h70, 8'h1d}; // CH=3 OP=0
cfg[2981] = { 1'b1, 8'haf, 8'hc6}; // CH=6 OP=3
cfg[2982] = { 1'b1, 8'h7a, 8'h1c}; // CH=5 OP=2
cfg[2983] = { 1'b0, 8'h5d, 8'hfc}; // CH=1 OP=3
cfg[2984] = { 1'b0, 8'h3e, 8'hb8}; // CH=2 OP=3
cfg[2985] = { 1'b1, 8'hc6, 8'h20}; // CH=5 OP=1
cfg[2986] = { 1'b0, 8'hc3, 8'h16}; // CH=3 OP=0
cfg[2987] = { 1'b1, 8'hc7, 8'h37}; // CH=6 OP=1
cfg[2988] = { 1'b0, 8'hc6, 8'h50}; // CH=2 OP=1
cfg[2989] = { 1'b0, 8'ha2, 8'ha6}; // CH=2 OP=0
cfg[2990] = { 1'b1, 8'h36, 8'hc3}; // CH=5 OP=1
cfg[2991] = { 1'b0, 8'hc9, 8'hc2}; // CH=1 OP=2
cfg[2992] = { 1'b0, 8'hcd, 8'h3c}; // CH=1 OP=3
cfg[2993] = { 1'b0, 8'h83, 8'h9a}; // CH=3 OP=0
cfg[2994] = { 1'b1, 8'hcd, 8'hd8}; // CH=4 OP=3
cfg[2995] = { 1'b1, 8'haf, 8'h9e}; // CH=6 OP=3
cfg[2996] = { 1'b0, 8'h57, 8'h61}; // CH=3 OP=1
cfg[2997] = { 1'b1, 8'h3b, 8'h28}; // CH=6 OP=2
cfg[2998] = { 1'b0, 8'h6c, 8'h33}; // CH=0 OP=3
cfg[2999] = { 1'b0, 8'h63, 8'ha3}; // CH=3 OP=0
cfg[3000] = { 1'b1, 8'h99, 8'hb5}; // CH=4 OP=2
cfg[3001] = { 1'b1, 8'h62, 8'h77}; // CH=5 OP=0
cfg[3002] = { 1'b0, 8'h70, 8'hb4}; // CH=0 OP=0
cfg[3003] = { 1'b0, 8'hcb, 8'hb3}; // CH=3 OP=2
cfg[3004] = { 1'b0, 8'h47, 8'h80}; // CH=3 OP=1
cfg[3005] = { 1'b0, 8'hd9, 8'h2f}; // CH=1 OP=2
cfg[3006] = { 1'b1, 8'ha2, 8'h86}; // CH=5 OP=0
cfg[3007] = { 1'b1, 8'hbc, 8'hc1}; // CH=3 OP=3
cfg[3008] = { 1'b0, 8'h5a, 8'hc2}; // CH=2 OP=2
cfg[3009] = { 1'b1, 8'hf8, 8'h8b}; // CH=3 OP=2
cfg[3010] = { 1'b1, 8'h92, 8'h24}; // CH=5 OP=0
cfg[3011] = { 1'b0, 8'h46, 8'hed}; // CH=2 OP=1
cfg[3012] = { 1'b0, 8'h94, 8'h5e}; // CH=0 OP=1
cfg[3013] = { 1'b1, 8'hba, 8'h29}; // CH=5 OP=2
cfg[3014] = { 1'b1, 8'h7e, 8'h70}; // CH=5 OP=3
cfg[3015] = { 1'b0, 8'ha3, 8'h49}; // CH=3 OP=0
cfg[3016] = { 1'b1, 8'hf0, 8'hec}; // CH=3 OP=0
cfg[3017] = { 1'b0, 8'h71, 8'ha8}; // CH=1 OP=0
cfg[3018] = { 1'b1, 8'hcb, 8'hd1}; // CH=6 OP=2
cfg[3019] = { 1'b0, 8'hc3, 8'h5c}; // CH=3 OP=0
cfg[3020] = { 1'b1, 8'he3, 8'h81}; // CH=6 OP=0
cfg[3021] = { 1'b0, 8'hd0, 8'h7}; // CH=0 OP=0
cfg[3022] = { 1'b0, 8'h58, 8'hbd}; // CH=0 OP=2
cfg[3023] = { 1'b1, 8'hc8, 8'hf}; // CH=3 OP=2
cfg[3024] = { 1'b0, 8'hed, 8'h28}; // CH=1 OP=3
cfg[3025] = { 1'b1, 8'hde, 8'hfe}; // CH=5 OP=3
cfg[3026] = { 1'b1, 8'h4f, 8'ha6}; // CH=6 OP=3
cfg[3027] = { 1'b0, 8'hd3, 8'h77}; // CH=3 OP=0
cfg[3028] = { 1'b0, 8'h76, 8'hde}; // CH=2 OP=1
cfg[3029] = { 1'b1, 8'hac, 8'hc1}; // CH=3 OP=3
cfg[3030] = { 1'b0, 8'hc0, 8'h91}; // CH=0 OP=0
cfg[3031] = { 1'b0, 8'h50, 8'h40}; // CH=0 OP=0
cfg[3032] = { 1'b0, 8'h78, 8'h4f}; // CH=0 OP=2
cfg[3033] = { 1'b0, 8'h3f, 8'h3d}; // CH=3 OP=3
cfg[3034] = { 1'b0, 8'h66, 8'h1b}; // CH=2 OP=1
cfg[3035] = { 1'b1, 8'hb1, 8'h6a}; // CH=4 OP=0
cfg[3036] = { 1'b0, 8'h84, 8'h84}; // CH=0 OP=1
cfg[3037] = { 1'b0, 8'hfa, 8'h62}; // CH=2 OP=2
cfg[3038] = { 1'b1, 8'ha7, 8'h23}; // CH=6 OP=1
cfg[3039] = { 1'b0, 8'hd0, 8'hb5}; // CH=0 OP=0
cfg[3040] = { 1'b0, 8'hee, 8'h75}; // CH=2 OP=3
cfg[3041] = { 1'b1, 8'h3e, 8'hf}; // CH=5 OP=3
cfg[3042] = { 1'b1, 8'hb6, 8'h5f}; // CH=5 OP=1
cfg[3043] = { 1'b0, 8'hf5, 8'h9c}; // CH=1 OP=1
cfg[3044] = { 1'b0, 8'h5c, 8'hb7}; // CH=0 OP=3
cfg[3045] = { 1'b1, 8'hf6, 8'h21}; // CH=5 OP=1
cfg[3046] = { 1'b1, 8'hd8, 8'h91}; // CH=3 OP=2
cfg[3047] = { 1'b0, 8'h32, 8'h8b}; // CH=2 OP=0
cfg[3048] = { 1'b0, 8'h52, 8'he0}; // CH=2 OP=0
cfg[3049] = { 1'b1, 8'h40, 8'hc}; // CH=3 OP=0
cfg[3050] = { 1'b0, 8'h7f, 8'h1c}; // CH=3 OP=3
cfg[3051] = { 1'b0, 8'h35, 8'h7b}; // CH=1 OP=1
cfg[3052] = { 1'b0, 8'hce, 8'h17}; // CH=2 OP=3
cfg[3053] = { 1'b1, 8'hef, 8'he8}; // CH=6 OP=3
cfg[3054] = { 1'b0, 8'h94, 8'hde}; // CH=0 OP=1
cfg[3055] = { 1'b1, 8'h9c, 8'hb6}; // CH=3 OP=3
cfg[3056] = { 1'b0, 8'hc8, 8'hc6}; // CH=0 OP=2
cfg[3057] = { 1'b1, 8'ha8, 8'h6a}; // CH=3 OP=2
cfg[3058] = { 1'b1, 8'hfe, 8'hbc}; // CH=5 OP=3
cfg[3059] = { 1'b0, 8'he0, 8'hfd}; // CH=0 OP=0
cfg[3060] = { 1'b0, 8'h30, 8'h7c}; // CH=0 OP=0
cfg[3061] = { 1'b1, 8'he0, 8'hb1}; // CH=3 OP=0
cfg[3062] = { 1'b0, 8'he1, 8'hdc}; // CH=1 OP=0
cfg[3063] = { 1'b0, 8'hc9, 8'h63}; // CH=1 OP=2
cfg[3064] = { 1'b1, 8'ha7, 8'hf7}; // CH=6 OP=1
cfg[3065] = { 1'b1, 8'h5d, 8'h1c}; // CH=4 OP=3
cfg[3066] = { 1'b0, 8'h56, 8'hcd}; // CH=2 OP=1
cfg[3067] = { 1'b0, 8'hfe, 8'h8e}; // CH=2 OP=3
cfg[3068] = { 1'b1, 8'hfc, 8'h4b}; // CH=3 OP=3
cfg[3069] = { 1'b1, 8'hdd, 8'h48}; // CH=4 OP=3
cfg[3070] = { 1'b1, 8'h75, 8'hc4}; // CH=4 OP=1
cfg[3071] = { 1'b0, 8'h52, 8'hbe}; // CH=2 OP=0
cfg[3072] = { 1'b1, 8'hb5, 8'h2c}; // CH=4 OP=1
cfg[3073] = { 1'b0, 8'had, 8'h89}; // CH=1 OP=3
cfg[3074] = { 1'b1, 8'hc9, 8'h7b}; // CH=4 OP=2
cfg[3075] = { 1'b0, 8'h96, 8'h9}; // CH=2 OP=1
cfg[3076] = { 1'b0, 8'h46, 8'h5f}; // CH=2 OP=1
cfg[3077] = { 1'b1, 8'hdc, 8'h5d}; // CH=3 OP=3
cfg[3078] = { 1'b0, 8'h63, 8'h5a}; // CH=3 OP=0
cfg[3079] = { 1'b0, 8'hf9, 8'h37}; // CH=1 OP=2
cfg[3080] = { 1'b0, 8'h32, 8'h44}; // CH=2 OP=0
cfg[3081] = { 1'b0, 8'h99, 8'h6d}; // CH=1 OP=2
cfg[3082] = { 1'b0, 8'hd8, 8'hd0}; // CH=0 OP=2
cfg[3083] = { 1'b1, 8'h75, 8'h99}; // CH=4 OP=1
cfg[3084] = { 1'b0, 8'h35, 8'h30}; // CH=1 OP=1
cfg[3085] = { 1'b1, 8'h84, 8'h76}; // CH=3 OP=1
cfg[3086] = { 1'b0, 8'hb6, 8'h52}; // CH=2 OP=1
cfg[3087] = { 1'b0, 8'haf, 8'h5d}; // CH=3 OP=3
cfg[3088] = { 1'b0, 8'hc6, 8'ha2}; // CH=2 OP=1
cfg[3089] = { 1'b0, 8'h9c, 8'hd4}; // CH=0 OP=3
cfg[3090] = { 1'b1, 8'h9f, 8'hd6}; // CH=6 OP=3
cfg[3091] = { 1'b0, 8'h48, 8'h6f}; // CH=0 OP=2
cfg[3092] = { 1'b0, 8'hbd, 8'hbc}; // CH=1 OP=3
cfg[3093] = { 1'b0, 8'hf2, 8'hec}; // CH=2 OP=0
cfg[3094] = { 1'b1, 8'h77, 8'h62}; // CH=6 OP=1
cfg[3095] = { 1'b1, 8'h95, 8'hb5}; // CH=4 OP=1
cfg[3096] = { 1'b0, 8'h96, 8'h6b}; // CH=2 OP=1
cfg[3097] = { 1'b1, 8'h3c, 8'h1a}; // CH=3 OP=3
cfg[3098] = { 1'b1, 8'hfe, 8'he0}; // CH=5 OP=3
cfg[3099] = { 1'b0, 8'h4e, 8'h7d}; // CH=2 OP=3
cfg[3100] = { 1'b0, 8'hbd, 8'h80}; // CH=1 OP=3
cfg[3101] = { 1'b1, 8'h79, 8'ha3}; // CH=4 OP=2
cfg[3102] = { 1'b1, 8'hbb, 8'hc2}; // CH=6 OP=2
cfg[3103] = { 1'b1, 8'h6c, 8'hb5}; // CH=3 OP=3
cfg[3104] = { 1'b1, 8'he9, 8'h2c}; // CH=4 OP=2
cfg[3105] = { 1'b0, 8'h8d, 8'hc1}; // CH=1 OP=3
cfg[3106] = { 1'b1, 8'h8f, 8'h57}; // CH=6 OP=3
cfg[3107] = { 1'b1, 8'h32, 8'h94}; // CH=5 OP=0
cfg[3108] = { 1'b0, 8'haa, 8'h92}; // CH=2 OP=2
cfg[3109] = { 1'b1, 8'hf8, 8'hc0}; // CH=3 OP=2
cfg[3110] = { 1'b1, 8'hb6, 8'h41}; // CH=5 OP=1
cfg[3111] = { 1'b0, 8'hbb, 8'he4}; // CH=3 OP=2
cfg[3112] = { 1'b1, 8'h7e, 8'h43}; // CH=5 OP=3
cfg[3113] = { 1'b0, 8'h33, 8'h8e}; // CH=3 OP=0
cfg[3114] = { 1'b0, 8'h5f, 8'h3b}; // CH=3 OP=3
cfg[3115] = { 1'b1, 8'hbf, 8'h9e}; // CH=6 OP=3
cfg[3116] = { 1'b1, 8'h4e, 8'h78}; // CH=5 OP=3
cfg[3117] = { 1'b1, 8'h80, 8'hc}; // CH=3 OP=0
cfg[3118] = { 1'b1, 8'h60, 8'h9e}; // CH=3 OP=0
cfg[3119] = { 1'b1, 8'hc1, 8'h23}; // CH=4 OP=0
cfg[3120] = { 1'b0, 8'h69, 8'hd9}; // CH=1 OP=2
cfg[3121] = { 1'b0, 8'h8a, 8'h95}; // CH=2 OP=2
cfg[3122] = { 1'b1, 8'h66, 8'h13}; // CH=5 OP=1
cfg[3123] = { 1'b1, 8'hae, 8'h46}; // CH=5 OP=3
cfg[3124] = { 1'b0, 8'hdf, 8'ha5}; // CH=3 OP=3
cfg[3125] = { 1'b0, 8'h9e, 8'hc5}; // CH=2 OP=3
cfg[3126] = { 1'b0, 8'hec, 8'h3d}; // CH=0 OP=3
cfg[3127] = { 1'b1, 8'h6d, 8'h49}; // CH=4 OP=3
cfg[3128] = { 1'b0, 8'h98, 8'he8}; // CH=0 OP=2
cfg[3129] = { 1'b0, 8'hbb, 8'h47}; // CH=3 OP=2
cfg[3130] = { 1'b1, 8'h95, 8'he7}; // CH=4 OP=1
cfg[3131] = { 1'b0, 8'h32, 8'h6b}; // CH=2 OP=0
cfg[3132] = { 1'b1, 8'h87, 8'h82}; // CH=6 OP=1
cfg[3133] = { 1'b1, 8'h46, 8'h30}; // CH=5 OP=1
cfg[3134] = { 1'b1, 8'he0, 8'hae}; // CH=3 OP=0
cfg[3135] = { 1'b1, 8'hcd, 8'h9a}; // CH=4 OP=3
cfg[3136] = { 1'b0, 8'hd5, 8'h7}; // CH=1 OP=1
cfg[3137] = { 1'b0, 8'h3d, 8'h9f}; // CH=1 OP=3
cfg[3138] = { 1'b1, 8'h66, 8'h5b}; // CH=5 OP=1
cfg[3139] = { 1'b0, 8'hf8, 8'hf0}; // CH=0 OP=2
cfg[3140] = { 1'b1, 8'h57, 8'h1a}; // CH=6 OP=1
cfg[3141] = { 1'b0, 8'hda, 8'hae}; // CH=2 OP=2
cfg[3142] = { 1'b0, 8'hd5, 8'hc6}; // CH=1 OP=1
cfg[3143] = { 1'b0, 8'h83, 8'hef}; // CH=3 OP=0
cfg[3144] = { 1'b0, 8'hb9, 8'h1a}; // CH=1 OP=2
cfg[3145] = { 1'b1, 8'h8e, 8'h25}; // CH=5 OP=3
cfg[3146] = { 1'b1, 8'hcb, 8'hc5}; // CH=6 OP=2
cfg[3147] = { 1'b1, 8'h31, 8'h20}; // CH=4 OP=0
cfg[3148] = { 1'b1, 8'h3d, 8'h10}; // CH=4 OP=3
cfg[3149] = { 1'b0, 8'hd3, 8'h81}; // CH=3 OP=0
cfg[3150] = { 1'b1, 8'h99, 8'h5b}; // CH=4 OP=2
cfg[3151] = { 1'b1, 8'h6e, 8'h5d}; // CH=5 OP=3
cfg[3152] = { 1'b1, 8'hf2, 8'h4c}; // CH=5 OP=0
cfg[3153] = { 1'b1, 8'h5c, 8'h67}; // CH=3 OP=3
cfg[3154] = { 1'b0, 8'hea, 8'h35}; // CH=2 OP=2
cfg[3155] = { 1'b1, 8'hb5, 8'hfa}; // CH=4 OP=1
cfg[3156] = { 1'b0, 8'he6, 8'h1a}; // CH=2 OP=1
cfg[3157] = { 1'b0, 8'h99, 8'h2a}; // CH=1 OP=2
cfg[3158] = { 1'b0, 8'hcf, 8'h4c}; // CH=3 OP=3
cfg[3159] = { 1'b1, 8'hb4, 8'h1f}; // CH=3 OP=1
cfg[3160] = { 1'b0, 8'h5f, 8'hb8}; // CH=3 OP=3
cfg[3161] = { 1'b1, 8'hda, 8'h26}; // CH=5 OP=2
cfg[3162] = { 1'b0, 8'h41, 8'hb9}; // CH=1 OP=0
cfg[3163] = { 1'b0, 8'h37, 8'h15}; // CH=3 OP=1
cfg[3164] = { 1'b0, 8'h58, 8'hff}; // CH=0 OP=2
cfg[3165] = { 1'b0, 8'h73, 8'h89}; // CH=3 OP=0
cfg[3166] = { 1'b0, 8'h9d, 8'h13}; // CH=1 OP=3
cfg[3167] = { 1'b1, 8'hf2, 8'hac}; // CH=5 OP=0
cfg[3168] = { 1'b1, 8'hc7, 8'h7b}; // CH=6 OP=1
cfg[3169] = { 1'b0, 8'hf8, 8'h30}; // CH=0 OP=2
cfg[3170] = { 1'b0, 8'h85, 8'h8f}; // CH=1 OP=1
cfg[3171] = { 1'b1, 8'h5f, 8'ha6}; // CH=6 OP=3
cfg[3172] = { 1'b1, 8'ha0, 8'h5f}; // CH=3 OP=0
cfg[3173] = { 1'b0, 8'hd7, 8'h75}; // CH=3 OP=1
cfg[3174] = { 1'b0, 8'hf0, 8'h74}; // CH=0 OP=0
cfg[3175] = { 1'b0, 8'h79, 8'h29}; // CH=1 OP=2
cfg[3176] = { 1'b1, 8'h8c, 8'hc3}; // CH=3 OP=3
cfg[3177] = { 1'b1, 8'h38, 8'h6d}; // CH=3 OP=2
cfg[3178] = { 1'b1, 8'hb3, 8'h62}; // CH=6 OP=0
cfg[3179] = { 1'b0, 8'he3, 8'h77}; // CH=3 OP=0
cfg[3180] = { 1'b0, 8'h73, 8'h43}; // CH=3 OP=0
cfg[3181] = { 1'b0, 8'h91, 8'h36}; // CH=1 OP=0
cfg[3182] = { 1'b0, 8'h32, 8'h78}; // CH=2 OP=0
cfg[3183] = { 1'b0, 8'h62, 8'hed}; // CH=2 OP=0
cfg[3184] = { 1'b1, 8'h8b, 8'hf2}; // CH=6 OP=2
cfg[3185] = { 1'b0, 8'h4e, 8'h50}; // CH=2 OP=3
cfg[3186] = { 1'b0, 8'hbb, 8'h4b}; // CH=3 OP=2
cfg[3187] = { 1'b0, 8'hea, 8'h38}; // CH=2 OP=2
cfg[3188] = { 1'b0, 8'hcd, 8'h95}; // CH=1 OP=3
cfg[3189] = { 1'b1, 8'h40, 8'hd8}; // CH=3 OP=0
cfg[3190] = { 1'b1, 8'h59, 8'hf}; // CH=4 OP=2
cfg[3191] = { 1'b0, 8'hd2, 8'h51}; // CH=2 OP=0
cfg[3192] = { 1'b0, 8'hbf, 8'hc7}; // CH=3 OP=3
cfg[3193] = { 1'b0, 8'h91, 8'hcf}; // CH=1 OP=0
cfg[3194] = { 1'b1, 8'hfb, 8'hac}; // CH=6 OP=2
cfg[3195] = { 1'b0, 8'hb6, 8'h5c}; // CH=2 OP=1
cfg[3196] = { 1'b1, 8'hd4, 8'h94}; // CH=3 OP=1
cfg[3197] = { 1'b1, 8'h69, 8'h81}; // CH=4 OP=2
cfg[3198] = { 1'b0, 8'h42, 8'h1a}; // CH=2 OP=0
cfg[3199] = { 1'b1, 8'h51, 8'he5}; // CH=4 OP=0
cfg[3200] = { 1'b0, 8'ha2, 8'h41}; // CH=2 OP=0
cfg[3201] = { 1'b0, 8'h69, 8'hd0}; // CH=1 OP=2
cfg[3202] = { 1'b0, 8'h38, 8'h68}; // CH=0 OP=2
cfg[3203] = { 1'b1, 8'hf9, 8'hf9}; // CH=4 OP=2
cfg[3204] = { 1'b0, 8'he5, 8'hfd}; // CH=1 OP=1
cfg[3205] = { 1'b0, 8'h9b, 8'h67}; // CH=3 OP=2
cfg[3206] = { 1'b1, 8'h70, 8'hfc}; // CH=3 OP=0
cfg[3207] = { 1'b0, 8'hd9, 8'h7d}; // CH=1 OP=2
cfg[3208] = { 1'b0, 8'h7d, 8'h97}; // CH=1 OP=3
cfg[3209] = { 1'b0, 8'hbd, 8'h6c}; // CH=1 OP=3
cfg[3210] = { 1'b0, 8'h8d, 8'h64}; // CH=1 OP=3
cfg[3211] = { 1'b1, 8'hf5, 8'h80}; // CH=4 OP=1
cfg[3212] = { 1'b1, 8'hef, 8'hbe}; // CH=6 OP=3
cfg[3213] = { 1'b1, 8'hec, 8'ha8}; // CH=3 OP=3
cfg[3214] = { 1'b0, 8'hec, 8'h8d}; // CH=0 OP=3
cfg[3215] = { 1'b1, 8'h98, 8'h28}; // CH=3 OP=2
cfg[3216] = { 1'b1, 8'h72, 8'h94}; // CH=5 OP=0
cfg[3217] = { 1'b0, 8'h8d, 8'h2b}; // CH=1 OP=3
cfg[3218] = { 1'b1, 8'hfa, 8'ha7}; // CH=5 OP=2
cfg[3219] = { 1'b1, 8'hb8, 8'h65}; // CH=3 OP=2
cfg[3220] = { 1'b0, 8'h38, 8'h80}; // CH=0 OP=2
cfg[3221] = { 1'b0, 8'hf6, 8'h2f}; // CH=2 OP=1
cfg[3222] = { 1'b1, 8'h9e, 8'hd8}; // CH=5 OP=3
cfg[3223] = { 1'b1, 8'hb0, 8'h8c}; // CH=3 OP=0
cfg[3224] = { 1'b0, 8'hd5, 8'h54}; // CH=1 OP=1
cfg[3225] = { 1'b1, 8'h57, 8'hec}; // CH=6 OP=1
cfg[3226] = { 1'b0, 8'h7f, 8'h5e}; // CH=3 OP=3
cfg[3227] = { 1'b0, 8'he6, 8'h70}; // CH=2 OP=1
cfg[3228] = { 1'b0, 8'hee, 8'h8c}; // CH=2 OP=3
cfg[3229] = { 1'b0, 8'h6e, 8'h7e}; // CH=2 OP=3
cfg[3230] = { 1'b0, 8'h9e, 8'h66}; // CH=2 OP=3
cfg[3231] = { 1'b1, 8'h76, 8'h3d}; // CH=5 OP=1
cfg[3232] = { 1'b1, 8'h75, 8'h1}; // CH=4 OP=1
cfg[3233] = { 1'b1, 8'hc9, 8'hab}; // CH=4 OP=2
cfg[3234] = { 1'b0, 8'hb5, 8'h6a}; // CH=1 OP=1
cfg[3235] = { 1'b1, 8'h3e, 8'hbe}; // CH=5 OP=3
cfg[3236] = { 1'b0, 8'h65, 8'h73}; // CH=1 OP=1
cfg[3237] = { 1'b0, 8'hf1, 8'h37}; // CH=1 OP=0
cfg[3238] = { 1'b0, 8'h6f, 8'hb3}; // CH=3 OP=3
cfg[3239] = { 1'b1, 8'hd6, 8'h67}; // CH=5 OP=1
cfg[3240] = { 1'b1, 8'h57, 8'h12}; // CH=6 OP=1
cfg[3241] = { 1'b0, 8'h5a, 8'h14}; // CH=2 OP=2
cfg[3242] = { 1'b1, 8'h9a, 8'hc5}; // CH=5 OP=2
cfg[3243] = { 1'b0, 8'h4f, 8'h70}; // CH=3 OP=3
cfg[3244] = { 1'b1, 8'h63, 8'h2e}; // CH=6 OP=0
cfg[3245] = { 1'b0, 8'h63, 8'h6c}; // CH=3 OP=0
cfg[3246] = { 1'b1, 8'h49, 8'hd1}; // CH=4 OP=2
cfg[3247] = { 1'b0, 8'h89, 8'hc2}; // CH=1 OP=2
cfg[3248] = { 1'b0, 8'hf0, 8'h61}; // CH=0 OP=0
cfg[3249] = { 1'b0, 8'h99, 8'h42}; // CH=1 OP=2
cfg[3250] = { 1'b1, 8'hf4, 8'h30}; // CH=3 OP=1
cfg[3251] = { 1'b0, 8'hf9, 8'hf5}; // CH=1 OP=2
cfg[3252] = { 1'b0, 8'h69, 8'h41}; // CH=1 OP=2
cfg[3253] = { 1'b1, 8'h98, 8'h6b}; // CH=3 OP=2
cfg[3254] = { 1'b1, 8'he0, 8'h97}; // CH=3 OP=0
cfg[3255] = { 1'b0, 8'h98, 8'hd6}; // CH=0 OP=2
cfg[3256] = { 1'b0, 8'hca, 8'h95}; // CH=2 OP=2
cfg[3257] = { 1'b1, 8'hd2, 8'h85}; // CH=5 OP=0
cfg[3258] = { 1'b1, 8'hee, 8'h88}; // CH=5 OP=3
cfg[3259] = { 1'b0, 8'h78, 8'he7}; // CH=0 OP=2
cfg[3260] = { 1'b1, 8'h72, 8'h13}; // CH=5 OP=0
cfg[3261] = { 1'b1, 8'hdb, 8'h55}; // CH=6 OP=2
cfg[3262] = { 1'b1, 8'h73, 8'hc0}; // CH=6 OP=0
cfg[3263] = { 1'b0, 8'h78, 8'h57}; // CH=0 OP=2
cfg[3264] = { 1'b0, 8'h4e, 8'h8d}; // CH=2 OP=3
cfg[3265] = { 1'b0, 8'he6, 8'h99}; // CH=2 OP=1
cfg[3266] = { 1'b0, 8'hb1, 8'h2e}; // CH=1 OP=0
cfg[3267] = { 1'b1, 8'h83, 8'hb3}; // CH=6 OP=0
cfg[3268] = { 1'b0, 8'h71, 8'h3c}; // CH=1 OP=0
cfg[3269] = { 1'b1, 8'h8f, 8'h23}; // CH=6 OP=3
cfg[3270] = { 1'b1, 8'ha3, 8'h3b}; // CH=6 OP=0
cfg[3271] = { 1'b1, 8'hf8, 8'h1c}; // CH=3 OP=2
cfg[3272] = { 1'b1, 8'hb8, 8'h17}; // CH=3 OP=2
cfg[3273] = { 1'b0, 8'h94, 8'h8f}; // CH=0 OP=1
cfg[3274] = { 1'b0, 8'he2, 8'h9c}; // CH=2 OP=0
cfg[3275] = { 1'b0, 8'hc9, 8'h35}; // CH=1 OP=2
cfg[3276] = { 1'b1, 8'h7a, 8'h63}; // CH=5 OP=2
cfg[3277] = { 1'b0, 8'hfd, 8'h16}; // CH=1 OP=3
cfg[3278] = { 1'b1, 8'h6f, 8'h52}; // CH=6 OP=3
cfg[3279] = { 1'b0, 8'hfe, 8'h76}; // CH=2 OP=3
cfg[3280] = { 1'b1, 8'ha1, 8'hb1}; // CH=4 OP=0
cfg[3281] = { 1'b1, 8'h99, 8'hcd}; // CH=4 OP=2
cfg[3282] = { 1'b0, 8'h51, 8'he5}; // CH=1 OP=0
cfg[3283] = { 1'b0, 8'h60, 8'h74}; // CH=0 OP=0
cfg[3284] = { 1'b1, 8'hfc, 8'h5c}; // CH=3 OP=3
cfg[3285] = { 1'b1, 8'h31, 8'hc7}; // CH=4 OP=0
cfg[3286] = { 1'b0, 8'h94, 8'hfc}; // CH=0 OP=1
cfg[3287] = { 1'b0, 8'hab, 8'ha4}; // CH=3 OP=2
cfg[3288] = { 1'b0, 8'hfd, 8'hab}; // CH=1 OP=3
cfg[3289] = { 1'b1, 8'h73, 8'h95}; // CH=6 OP=0
cfg[3290] = { 1'b1, 8'h9f, 8'hdb}; // CH=6 OP=3
cfg[3291] = { 1'b0, 8'h38, 8'hf2}; // CH=0 OP=2
cfg[3292] = { 1'b0, 8'h8a, 8'hd7}; // CH=2 OP=2
cfg[3293] = { 1'b0, 8'hea, 8'h4b}; // CH=2 OP=2
cfg[3294] = { 1'b1, 8'he7, 8'ha8}; // CH=6 OP=1
cfg[3295] = { 1'b1, 8'h57, 8'h6f}; // CH=6 OP=1
cfg[3296] = { 1'b1, 8'hea, 8'had}; // CH=5 OP=2
cfg[3297] = { 1'b1, 8'h7a, 8'h58}; // CH=5 OP=2
cfg[3298] = { 1'b1, 8'h79, 8'h55}; // CH=4 OP=2
cfg[3299] = { 1'b0, 8'h76, 8'hc9}; // CH=2 OP=1
cfg[3300] = { 1'b1, 8'hdf, 8'hed}; // CH=6 OP=3
cfg[3301] = { 1'b0, 8'hb6, 8'hc3}; // CH=2 OP=1
cfg[3302] = { 1'b0, 8'hc2, 8'h46}; // CH=2 OP=0
cfg[3303] = { 1'b1, 8'ha9, 8'haa}; // CH=4 OP=2
cfg[3304] = { 1'b0, 8'hc2, 8'h19}; // CH=2 OP=0
cfg[3305] = { 1'b0, 8'h6f, 8'h84}; // CH=3 OP=3
cfg[3306] = { 1'b0, 8'hc7, 8'h93}; // CH=3 OP=1
cfg[3307] = { 1'b0, 8'ha9, 8'h4e}; // CH=1 OP=2
cfg[3308] = { 1'b1, 8'hca, 8'he5}; // CH=5 OP=2
cfg[3309] = { 1'b1, 8'he4, 8'h35}; // CH=3 OP=1
cfg[3310] = { 1'b0, 8'ha7, 8'h83}; // CH=3 OP=1
cfg[3311] = { 1'b1, 8'hed, 8'h5b}; // CH=4 OP=3
cfg[3312] = { 1'b1, 8'hc7, 8'h1d}; // CH=6 OP=1
cfg[3313] = { 1'b1, 8'h89, 8'h2e}; // CH=4 OP=2
cfg[3314] = { 1'b1, 8'hf8, 8'hb2}; // CH=3 OP=2
cfg[3315] = { 1'b1, 8'hbf, 8'h45}; // CH=6 OP=3
cfg[3316] = { 1'b1, 8'hdb, 8'h94}; // CH=6 OP=2
cfg[3317] = { 1'b0, 8'hc1, 8'h33}; // CH=1 OP=0
cfg[3318] = { 1'b0, 8'h94, 8'hfd}; // CH=0 OP=1
cfg[3319] = { 1'b1, 8'h46, 8'he1}; // CH=5 OP=1
cfg[3320] = { 1'b0, 8'haf, 8'h89}; // CH=3 OP=3
cfg[3321] = { 1'b1, 8'h42, 8'h76}; // CH=5 OP=0
cfg[3322] = { 1'b1, 8'h31, 8'h2f}; // CH=4 OP=0
cfg[3323] = { 1'b1, 8'h94, 8'h92}; // CH=3 OP=1
cfg[3324] = { 1'b1, 8'hae, 8'h8a}; // CH=5 OP=3
cfg[3325] = { 1'b1, 8'hf7, 8'h49}; // CH=6 OP=1
cfg[3326] = { 1'b1, 8'hea, 8'h25}; // CH=5 OP=2
cfg[3327] = { 1'b0, 8'hfc, 8'he6}; // CH=0 OP=3
cfg[3328] = { 1'b1, 8'h43, 8'h7a}; // CH=6 OP=0
cfg[3329] = { 1'b1, 8'h84, 8'hc0}; // CH=3 OP=1
cfg[3330] = { 1'b0, 8'hfa, 8'h32}; // CH=2 OP=2
cfg[3331] = { 1'b0, 8'h94, 8'h74}; // CH=0 OP=1
cfg[3332] = { 1'b0, 8'hc5, 8'h7e}; // CH=1 OP=1
cfg[3333] = { 1'b1, 8'h59, 8'h10}; // CH=4 OP=2
cfg[3334] = { 1'b1, 8'h7c, 8'h9b}; // CH=3 OP=3
cfg[3335] = { 1'b0, 8'h65, 8'hff}; // CH=1 OP=1
cfg[3336] = { 1'b1, 8'h81, 8'he9}; // CH=4 OP=0
cfg[3337] = { 1'b1, 8'h9a, 8'he5}; // CH=5 OP=2
cfg[3338] = { 1'b1, 8'h95, 8'h28}; // CH=4 OP=1
cfg[3339] = { 1'b0, 8'h9a, 8'h35}; // CH=2 OP=2
cfg[3340] = { 1'b1, 8'hdb, 8'h14}; // CH=6 OP=2
cfg[3341] = { 1'b0, 8'h59, 8'hde}; // CH=1 OP=2
cfg[3342] = { 1'b1, 8'h6a, 8'hf6}; // CH=5 OP=2
cfg[3343] = { 1'b0, 8'hce, 8'h1d}; // CH=2 OP=3
cfg[3344] = { 1'b1, 8'hcd, 8'he9}; // CH=4 OP=3
cfg[3345] = { 1'b0, 8'hb6, 8'hf3}; // CH=2 OP=1
cfg[3346] = { 1'b1, 8'h9b, 8'he2}; // CH=6 OP=2
cfg[3347] = { 1'b1, 8'hc3, 8'h4c}; // CH=6 OP=0
cfg[3348] = { 1'b1, 8'hf8, 8'h76}; // CH=3 OP=2
cfg[3349] = { 1'b0, 8'h5f, 8'h10}; // CH=3 OP=3
cfg[3350] = { 1'b0, 8'h3a, 8'h34}; // CH=2 OP=2
cfg[3351] = { 1'b0, 8'h94, 8'h13}; // CH=0 OP=1
cfg[3352] = { 1'b1, 8'hfe, 8'h9}; // CH=5 OP=3
cfg[3353] = { 1'b0, 8'h86, 8'h26}; // CH=2 OP=1
cfg[3354] = { 1'b1, 8'h53, 8'hec}; // CH=6 OP=0
cfg[3355] = { 1'b1, 8'h3c, 8'hdf}; // CH=3 OP=3
cfg[3356] = { 1'b0, 8'h55, 8'ha4}; // CH=1 OP=1
cfg[3357] = { 1'b0, 8'h84, 8'h67}; // CH=0 OP=1
cfg[3358] = { 1'b1, 8'h94, 8'hcd}; // CH=3 OP=1
cfg[3359] = { 1'b0, 8'hc8, 8'ha9}; // CH=0 OP=2
cfg[3360] = { 1'b0, 8'hdb, 8'h2e}; // CH=3 OP=2
cfg[3361] = { 1'b0, 8'he4, 8'h1f}; // CH=0 OP=1
cfg[3362] = { 1'b0, 8'h8d, 8'hd7}; // CH=1 OP=3
cfg[3363] = { 1'b1, 8'h7a, 8'hc9}; // CH=5 OP=2
cfg[3364] = { 1'b0, 8'h59, 8'h86}; // CH=1 OP=2
cfg[3365] = { 1'b1, 8'h5d, 8'hc2}; // CH=4 OP=3
cfg[3366] = { 1'b0, 8'hc4, 8'h29}; // CH=0 OP=1
cfg[3367] = { 1'b0, 8'he9, 8'had}; // CH=1 OP=2
cfg[3368] = { 1'b1, 8'h93, 8'he1}; // CH=6 OP=0
cfg[3369] = { 1'b0, 8'hc1, 8'hda}; // CH=1 OP=0
cfg[3370] = { 1'b1, 8'he0, 8'h66}; // CH=3 OP=0
cfg[3371] = { 1'b0, 8'hb8, 8'hf1}; // CH=0 OP=2
cfg[3372] = { 1'b0, 8'h9e, 8'h7e}; // CH=2 OP=3
cfg[3373] = { 1'b0, 8'h52, 8'hc6}; // CH=2 OP=0
cfg[3374] = { 1'b1, 8'h6d, 8'he7}; // CH=4 OP=3
cfg[3375] = { 1'b1, 8'h97, 8'hff}; // CH=6 OP=1
cfg[3376] = { 1'b1, 8'h44, 8'h1b}; // CH=3 OP=1
cfg[3377] = { 1'b1, 8'h86, 8'h5}; // CH=5 OP=1
cfg[3378] = { 1'b0, 8'h90, 8'h98}; // CH=0 OP=0
cfg[3379] = { 1'b0, 8'h75, 8'h59}; // CH=1 OP=1
cfg[3380] = { 1'b1, 8'h3f, 8'h39}; // CH=6 OP=3
cfg[3381] = { 1'b0, 8'h56, 8'hf1}; // CH=2 OP=1
cfg[3382] = { 1'b1, 8'h4f, 8'hb2}; // CH=6 OP=3
cfg[3383] = { 1'b1, 8'ha1, 8'hd6}; // CH=4 OP=0
cfg[3384] = { 1'b0, 8'hbc, 8'hbd}; // CH=0 OP=3
cfg[3385] = { 1'b1, 8'hd8, 8'hcb}; // CH=3 OP=2
cfg[3386] = { 1'b0, 8'hdd, 8'h90}; // CH=1 OP=3
cfg[3387] = { 1'b0, 8'h75, 8'h36}; // CH=1 OP=1
cfg[3388] = { 1'b0, 8'hce, 8'hb7}; // CH=2 OP=3
cfg[3389] = { 1'b1, 8'hb5, 8'h9e}; // CH=4 OP=1
cfg[3390] = { 1'b0, 8'hc9, 8'hf9}; // CH=1 OP=2
cfg[3391] = { 1'b0, 8'h7b, 8'h0}; // CH=3 OP=2
cfg[3392] = { 1'b1, 8'h51, 8'hcd}; // CH=4 OP=0
cfg[3393] = { 1'b0, 8'hcb, 8'h19}; // CH=3 OP=2
cfg[3394] = { 1'b1, 8'h70, 8'hcb}; // CH=3 OP=0
cfg[3395] = { 1'b0, 8'h5a, 8'ha3}; // CH=2 OP=2
cfg[3396] = { 1'b0, 8'hca, 8'h80}; // CH=2 OP=2
cfg[3397] = { 1'b0, 8'hca, 8'hf5}; // CH=2 OP=2
cfg[3398] = { 1'b1, 8'h40, 8'hc3}; // CH=3 OP=0
cfg[3399] = { 1'b1, 8'hf5, 8'hcb}; // CH=4 OP=1
cfg[3400] = { 1'b1, 8'hbe, 8'hc4}; // CH=5 OP=3
cfg[3401] = { 1'b0, 8'h39, 8'hc4}; // CH=1 OP=2
cfg[3402] = { 1'b1, 8'h8a, 8'h91}; // CH=5 OP=2
cfg[3403] = { 1'b0, 8'h99, 8'haa}; // CH=1 OP=2
cfg[3404] = { 1'b1, 8'h65, 8'hed}; // CH=4 OP=1
cfg[3405] = { 1'b1, 8'hda, 8'hfb}; // CH=5 OP=2
cfg[3406] = { 1'b1, 8'ha4, 8'h89}; // CH=3 OP=1
cfg[3407] = { 1'b0, 8'h6f, 8'h7e}; // CH=3 OP=3
cfg[3408] = { 1'b1, 8'haf, 8'h42}; // CH=6 OP=3
cfg[3409] = { 1'b1, 8'ha4, 8'hd}; // CH=3 OP=1
cfg[3410] = { 1'b0, 8'h62, 8'hd1}; // CH=2 OP=0
cfg[3411] = { 1'b0, 8'h9b, 8'h95}; // CH=3 OP=2
cfg[3412] = { 1'b0, 8'hfa, 8'h26}; // CH=2 OP=2
cfg[3413] = { 1'b0, 8'hbe, 8'hbf}; // CH=2 OP=3
cfg[3414] = { 1'b0, 8'hb9, 8'h88}; // CH=1 OP=2
cfg[3415] = { 1'b0, 8'h53, 8'h62}; // CH=3 OP=0
cfg[3416] = { 1'b1, 8'hc1, 8'h7}; // CH=4 OP=0
cfg[3417] = { 1'b0, 8'hba, 8'h76}; // CH=2 OP=2
cfg[3418] = { 1'b0, 8'hdd, 8'h25}; // CH=1 OP=3
cfg[3419] = { 1'b1, 8'ha0, 8'hc9}; // CH=3 OP=0
cfg[3420] = { 1'b0, 8'hce, 8'h2b}; // CH=2 OP=3
cfg[3421] = { 1'b1, 8'h84, 8'hc6}; // CH=3 OP=1
cfg[3422] = { 1'b1, 8'h7e, 8'heb}; // CH=5 OP=3
cfg[3423] = { 1'b1, 8'h87, 8'haa}; // CH=6 OP=1
cfg[3424] = { 1'b1, 8'h57, 8'hce}; // CH=6 OP=1
cfg[3425] = { 1'b1, 8'haa, 8'h72}; // CH=5 OP=2
cfg[3426] = { 1'b0, 8'h6b, 8'h79}; // CH=3 OP=2
cfg[3427] = { 1'b0, 8'h5a, 8'hef}; // CH=2 OP=2
cfg[3428] = { 1'b0, 8'hdd, 8'h3}; // CH=1 OP=3
cfg[3429] = { 1'b1, 8'h31, 8'ha3}; // CH=4 OP=0
cfg[3430] = { 1'b0, 8'hce, 8'h71}; // CH=2 OP=3
cfg[3431] = { 1'b0, 8'hba, 8'h29}; // CH=2 OP=2
cfg[3432] = { 1'b0, 8'h64, 8'h9}; // CH=0 OP=1
cfg[3433] = { 1'b0, 8'h33, 8'ha6}; // CH=3 OP=0
cfg[3434] = { 1'b0, 8'h7e, 8'hfd}; // CH=2 OP=3
cfg[3435] = { 1'b1, 8'hf8, 8'hde}; // CH=3 OP=2
cfg[3436] = { 1'b0, 8'he7, 8'hc3}; // CH=3 OP=1
cfg[3437] = { 1'b0, 8'hfc, 8'h1d}; // CH=0 OP=3
cfg[3438] = { 1'b1, 8'hd9, 8'hfb}; // CH=4 OP=2
cfg[3439] = { 1'b0, 8'he2, 8'h2c}; // CH=2 OP=0
cfg[3440] = { 1'b1, 8'hb0, 8'h47}; // CH=3 OP=0
cfg[3441] = { 1'b1, 8'h6a, 8'h70}; // CH=5 OP=2
cfg[3442] = { 1'b0, 8'hcf, 8'h79}; // CH=3 OP=3
cfg[3443] = { 1'b0, 8'hc2, 8'h20}; // CH=2 OP=0
cfg[3444] = { 1'b1, 8'h40, 8'h30}; // CH=3 OP=0
cfg[3445] = { 1'b1, 8'h38, 8'he}; // CH=3 OP=2
cfg[3446] = { 1'b1, 8'hef, 8'hd1}; // CH=6 OP=3
cfg[3447] = { 1'b0, 8'hea, 8'h4a}; // CH=2 OP=2
cfg[3448] = { 1'b1, 8'hd7, 8'h28}; // CH=6 OP=1
cfg[3449] = { 1'b0, 8'h88, 8'h5d}; // CH=0 OP=2
cfg[3450] = { 1'b1, 8'hf2, 8'hce}; // CH=5 OP=0
cfg[3451] = { 1'b1, 8'hc1, 8'h47}; // CH=4 OP=0
cfg[3452] = { 1'b1, 8'hc3, 8'h67}; // CH=6 OP=0
cfg[3453] = { 1'b1, 8'hf3, 8'h85}; // CH=6 OP=0
cfg[3454] = { 1'b0, 8'h68, 8'h4a}; // CH=0 OP=2
cfg[3455] = { 1'b1, 8'h88, 8'hd3}; // CH=3 OP=2
cfg[3456] = { 1'b1, 8'ha4, 8'hc2}; // CH=3 OP=1
cfg[3457] = { 1'b1, 8'h9a, 8'hac}; // CH=5 OP=2
cfg[3458] = { 1'b0, 8'h71, 8'hc3}; // CH=1 OP=0
cfg[3459] = { 1'b0, 8'hf9, 8'h20}; // CH=1 OP=2
cfg[3460] = { 1'b1, 8'hec, 8'hee}; // CH=3 OP=3
cfg[3461] = { 1'b1, 8'had, 8'h36}; // CH=4 OP=3
cfg[3462] = { 1'b0, 8'h71, 8'h9d}; // CH=1 OP=0
cfg[3463] = { 1'b0, 8'h64, 8'h22}; // CH=0 OP=1
cfg[3464] = { 1'b0, 8'h66, 8'h6c}; // CH=2 OP=1
cfg[3465] = { 1'b0, 8'h3a, 8'h8e}; // CH=2 OP=2
cfg[3466] = { 1'b1, 8'hfc, 8'hbf}; // CH=3 OP=3
cfg[3467] = { 1'b1, 8'ha9, 8'h3a}; // CH=4 OP=2
cfg[3468] = { 1'b1, 8'h6c, 8'hde}; // CH=3 OP=3
cfg[3469] = { 1'b1, 8'h8c, 8'hfa}; // CH=3 OP=3
cfg[3470] = { 1'b0, 8'h7b, 8'hd4}; // CH=3 OP=2
cfg[3471] = { 1'b0, 8'hb1, 8'h25}; // CH=1 OP=0
cfg[3472] = { 1'b0, 8'h4e, 8'ha3}; // CH=2 OP=3
cfg[3473] = { 1'b1, 8'h71, 8'h11}; // CH=4 OP=0
cfg[3474] = { 1'b1, 8'hdd, 8'haf}; // CH=4 OP=3
cfg[3475] = { 1'b0, 8'h6b, 8'hb6}; // CH=3 OP=2
cfg[3476] = { 1'b0, 8'h44, 8'h45}; // CH=0 OP=1
cfg[3477] = { 1'b0, 8'hed, 8'h65}; // CH=1 OP=3
cfg[3478] = { 1'b0, 8'h59, 8'h43}; // CH=1 OP=2
cfg[3479] = { 1'b1, 8'he6, 8'h3e}; // CH=5 OP=1
cfg[3480] = { 1'b1, 8'h61, 8'h12}; // CH=4 OP=0
cfg[3481] = { 1'b0, 8'hb4, 8'h37}; // CH=0 OP=1
cfg[3482] = { 1'b0, 8'hf7, 8'h60}; // CH=3 OP=1
cfg[3483] = { 1'b0, 8'h9e, 8'hd1}; // CH=2 OP=3
cfg[3484] = { 1'b1, 8'hac, 8'haf}; // CH=3 OP=3
cfg[3485] = { 1'b1, 8'hf4, 8'h1a}; // CH=3 OP=1
cfg[3486] = { 1'b0, 8'h39, 8'h45}; // CH=1 OP=2
cfg[3487] = { 1'b1, 8'h55, 8'haa}; // CH=4 OP=1
cfg[3488] = { 1'b1, 8'hda, 8'h80}; // CH=5 OP=2
cfg[3489] = { 1'b1, 8'h97, 8'h66}; // CH=6 OP=1
cfg[3490] = { 1'b1, 8'h79, 8'hc7}; // CH=4 OP=2
cfg[3491] = { 1'b0, 8'h4f, 8'hd9}; // CH=3 OP=3
cfg[3492] = { 1'b1, 8'h3b, 8'h24}; // CH=6 OP=2
cfg[3493] = { 1'b1, 8'hd6, 8'hc3}; // CH=5 OP=1
cfg[3494] = { 1'b0, 8'hd4, 8'h6f}; // CH=0 OP=1
cfg[3495] = { 1'b0, 8'h9d, 8'hbe}; // CH=1 OP=3
cfg[3496] = { 1'b1, 8'hc3, 8'hc3}; // CH=6 OP=0
cfg[3497] = { 1'b0, 8'h43, 8'hb1}; // CH=3 OP=0
cfg[3498] = { 1'b0, 8'ha9, 8'hdc}; // CH=1 OP=2
cfg[3499] = { 1'b0, 8'h70, 8'h1a}; // CH=0 OP=0
cfg[3500] = { 1'b1, 8'h49, 8'h8e}; // CH=4 OP=2
cfg[3501] = { 1'b1, 8'h83, 8'hdd}; // CH=6 OP=0
cfg[3502] = { 1'b1, 8'h8e, 8'h18}; // CH=5 OP=3
cfg[3503] = { 1'b0, 8'h48, 8'hef}; // CH=0 OP=2
cfg[3504] = { 1'b0, 8'hf6, 8'h17}; // CH=2 OP=1
cfg[3505] = { 1'b1, 8'h93, 8'h36}; // CH=6 OP=0
cfg[3506] = { 1'b1, 8'h56, 8'hf9}; // CH=5 OP=1
cfg[3507] = { 1'b1, 8'h9a, 8'haa}; // CH=5 OP=2
cfg[3508] = { 1'b0, 8'h43, 8'h87}; // CH=3 OP=0
cfg[3509] = { 1'b0, 8'hb4, 8'ha1}; // CH=0 OP=1
cfg[3510] = { 1'b1, 8'hfd, 8'h2f}; // CH=4 OP=3
cfg[3511] = { 1'b0, 8'h80, 8'hd}; // CH=0 OP=0
cfg[3512] = { 1'b0, 8'h56, 8'h25}; // CH=2 OP=1
cfg[3513] = { 1'b0, 8'h73, 8'h2b}; // CH=3 OP=0
cfg[3514] = { 1'b0, 8'ha9, 8'h1}; // CH=1 OP=2
cfg[3515] = { 1'b1, 8'ha2, 8'ha4}; // CH=5 OP=0
cfg[3516] = { 1'b0, 8'h4d, 8'h69}; // CH=1 OP=3
cfg[3517] = { 1'b0, 8'hd4, 8'h2b}; // CH=0 OP=1
cfg[3518] = { 1'b1, 8'h75, 8'h81}; // CH=4 OP=1
cfg[3519] = { 1'b1, 8'ha4, 8'he5}; // CH=3 OP=1
cfg[3520] = { 1'b1, 8'hb1, 8'h83}; // CH=4 OP=0
cfg[3521] = { 1'b1, 8'hd7, 8'h81}; // CH=6 OP=1
cfg[3522] = { 1'b0, 8'heb, 8'ha2}; // CH=3 OP=2
cfg[3523] = { 1'b0, 8'h79, 8'h54}; // CH=1 OP=2
cfg[3524] = { 1'b1, 8'h38, 8'h18}; // CH=3 OP=2
cfg[3525] = { 1'b0, 8'hca, 8'hc5}; // CH=2 OP=2
cfg[3526] = { 1'b1, 8'hf6, 8'h12}; // CH=5 OP=1
cfg[3527] = { 1'b1, 8'h66, 8'he6}; // CH=5 OP=1
cfg[3528] = { 1'b0, 8'h89, 8'h5b}; // CH=1 OP=2
cfg[3529] = { 1'b1, 8'haa, 8'hff}; // CH=5 OP=2
cfg[3530] = { 1'b1, 8'h4c, 8'hb1}; // CH=3 OP=3
cfg[3531] = { 1'b0, 8'hfc, 8'h88}; // CH=0 OP=3
cfg[3532] = { 1'b0, 8'hb3, 8'h73}; // CH=3 OP=0
cfg[3533] = { 1'b0, 8'hb0, 8'h7c}; // CH=0 OP=0
cfg[3534] = { 1'b0, 8'he8, 8'h9e}; // CH=0 OP=2
cfg[3535] = { 1'b0, 8'hb3, 8'h63}; // CH=3 OP=0
cfg[3536] = { 1'b0, 8'ha9, 8'h75}; // CH=1 OP=2
cfg[3537] = { 1'b1, 8'ha7, 8'h5b}; // CH=6 OP=1
cfg[3538] = { 1'b0, 8'h5f, 8'h99}; // CH=3 OP=3
cfg[3539] = { 1'b0, 8'h9a, 8'h43}; // CH=2 OP=2
cfg[3540] = { 1'b1, 8'h56, 8'h8f}; // CH=5 OP=1
cfg[3541] = { 1'b1, 8'hb5, 8'h8b}; // CH=4 OP=1
cfg[3542] = { 1'b0, 8'h68, 8'h8e}; // CH=0 OP=2
cfg[3543] = { 1'b1, 8'h8f, 8'ha}; // CH=6 OP=3
cfg[3544] = { 1'b0, 8'hee, 8'h0}; // CH=2 OP=3
cfg[3545] = { 1'b0, 8'h72, 8'hb3}; // CH=2 OP=0
cfg[3546] = { 1'b1, 8'h47, 8'h5d}; // CH=6 OP=1
cfg[3547] = { 1'b1, 8'hee, 8'h6c}; // CH=5 OP=3
cfg[3548] = { 1'b1, 8'h4d, 8'h5}; // CH=4 OP=3
cfg[3549] = { 1'b1, 8'he7, 8'h49}; // CH=6 OP=1
cfg[3550] = { 1'b0, 8'h3e, 8'hd8}; // CH=2 OP=3
cfg[3551] = { 1'b1, 8'hf3, 8'h64}; // CH=6 OP=0
cfg[3552] = { 1'b0, 8'h5b, 8'hf2}; // CH=3 OP=2
cfg[3553] = { 1'b1, 8'h73, 8'hfc}; // CH=6 OP=0
cfg[3554] = { 1'b0, 8'h73, 8'ha4}; // CH=3 OP=0
cfg[3555] = { 1'b0, 8'hde, 8'hb0}; // CH=2 OP=3
cfg[3556] = { 1'b0, 8'hf0, 8'h84}; // CH=0 OP=0
cfg[3557] = { 1'b0, 8'hf6, 8'ha2}; // CH=2 OP=1
cfg[3558] = { 1'b1, 8'h3f, 8'hec}; // CH=6 OP=3
cfg[3559] = { 1'b1, 8'h87, 8'h9c}; // CH=6 OP=1
cfg[3560] = { 1'b0, 8'h7a, 8'h7b}; // CH=2 OP=2
cfg[3561] = { 1'b0, 8'hd5, 8'h6d}; // CH=1 OP=1
cfg[3562] = { 1'b1, 8'h48, 8'h69}; // CH=3 OP=2
cfg[3563] = { 1'b1, 8'hbb, 8'he}; // CH=6 OP=2
cfg[3564] = { 1'b0, 8'he2, 8'hbe}; // CH=2 OP=0
cfg[3565] = { 1'b0, 8'h66, 8'hf0}; // CH=2 OP=1
cfg[3566] = { 1'b0, 8'h57, 8'hff}; // CH=3 OP=1
cfg[3567] = { 1'b0, 8'h4d, 8'ha2}; // CH=1 OP=3
cfg[3568] = { 1'b1, 8'h8c, 8'h8e}; // CH=3 OP=3
cfg[3569] = { 1'b0, 8'ha3, 8'h2a}; // CH=3 OP=0
cfg[3570] = { 1'b1, 8'hdb, 8'h66}; // CH=6 OP=2
cfg[3571] = { 1'b0, 8'hb0, 8'h8c}; // CH=0 OP=0
cfg[3572] = { 1'b1, 8'hf8, 8'hf6}; // CH=3 OP=2
cfg[3573] = { 1'b1, 8'hb4, 8'h4}; // CH=3 OP=1
cfg[3574] = { 1'b1, 8'h96, 8'hc2}; // CH=5 OP=1
cfg[3575] = { 1'b1, 8'hfd, 8'hb3}; // CH=4 OP=3
cfg[3576] = { 1'b1, 8'h54, 8'hb2}; // CH=3 OP=1
cfg[3577] = { 1'b1, 8'ha1, 8'h54}; // CH=4 OP=0
cfg[3578] = { 1'b1, 8'h43, 8'he2}; // CH=6 OP=0
cfg[3579] = { 1'b1, 8'ha5, 8'hd0}; // CH=4 OP=1
cfg[3580] = { 1'b1, 8'h80, 8'hef}; // CH=3 OP=0
cfg[3581] = { 1'b0, 8'h31, 8'h7c}; // CH=1 OP=0
cfg[3582] = { 1'b1, 8'h66, 8'h72}; // CH=5 OP=1
cfg[3583] = { 1'b0, 8'hfb, 8'hdd}; // CH=3 OP=2
cfg[3584] = { 1'b0, 8'h87, 8'h74}; // CH=3 OP=1
cfg[3585] = { 1'b1, 8'h9e, 8'h71}; // CH=5 OP=3
cfg[3586] = { 1'b1, 8'hf2, 8'h6}; // CH=5 OP=0
cfg[3587] = { 1'b0, 8'hd5, 8'h6f}; // CH=1 OP=1
cfg[3588] = { 1'b1, 8'he2, 8'hb2}; // CH=5 OP=0
cfg[3589] = { 1'b1, 8'h55, 8'h57}; // CH=4 OP=1
cfg[3590] = { 1'b1, 8'h6d, 8'hd8}; // CH=4 OP=3
cfg[3591] = { 1'b1, 8'h57, 8'h9}; // CH=6 OP=1
cfg[3592] = { 1'b1, 8'hbd, 8'h32}; // CH=4 OP=3
cfg[3593] = { 1'b1, 8'hb9, 8'h10}; // CH=4 OP=2
cfg[3594] = { 1'b1, 8'h40, 8'h84}; // CH=3 OP=0
cfg[3595] = { 1'b1, 8'h6e, 8'hf5}; // CH=5 OP=3
cfg[3596] = { 1'b1, 8'h74, 8'hba}; // CH=3 OP=1
cfg[3597] = { 1'b1, 8'he3, 8'h20}; // CH=6 OP=0
cfg[3598] = { 1'b0, 8'h96, 8'hb3}; // CH=2 OP=1
cfg[3599] = { 1'b0, 8'hed, 8'h16}; // CH=1 OP=3
cfg[3600] = { 1'b0, 8'hc5, 8'h69}; // CH=1 OP=1
cfg[3601] = { 1'b1, 8'hce, 8'h38}; // CH=5 OP=3
cfg[3602] = { 1'b0, 8'hfa, 8'h79}; // CH=2 OP=2
cfg[3603] = { 1'b0, 8'hb3, 8'h11}; // CH=3 OP=0
cfg[3604] = { 1'b0, 8'hf3, 8'h95}; // CH=3 OP=0
cfg[3605] = { 1'b1, 8'h61, 8'h8a}; // CH=4 OP=0
cfg[3606] = { 1'b0, 8'hd6, 8'h44}; // CH=2 OP=1
cfg[3607] = { 1'b1, 8'hb9, 8'h64}; // CH=4 OP=2
cfg[3608] = { 1'b0, 8'h4f, 8'h17}; // CH=3 OP=3
cfg[3609] = { 1'b0, 8'h3d, 8'h2d}; // CH=1 OP=3
cfg[3610] = { 1'b0, 8'ha0, 8'h97}; // CH=0 OP=0
cfg[3611] = { 1'b1, 8'hdc, 8'hd1}; // CH=3 OP=3
cfg[3612] = { 1'b1, 8'hd6, 8'hd2}; // CH=5 OP=1
cfg[3613] = { 1'b1, 8'h89, 8'he3}; // CH=4 OP=2
cfg[3614] = { 1'b1, 8'h7c, 8'h78}; // CH=3 OP=3
cfg[3615] = { 1'b0, 8'hde, 8'h2}; // CH=2 OP=3
cfg[3616] = { 1'b0, 8'hb4, 8'h46}; // CH=0 OP=1
cfg[3617] = { 1'b0, 8'h6d, 8'haa}; // CH=1 OP=3
cfg[3618] = { 1'b0, 8'hbd, 8'hc1}; // CH=1 OP=3
cfg[3619] = { 1'b0, 8'hfa, 8'hee}; // CH=2 OP=2
cfg[3620] = { 1'b1, 8'hfc, 8'h85}; // CH=3 OP=3
cfg[3621] = { 1'b1, 8'hcd, 8'h55}; // CH=4 OP=3
cfg[3622] = { 1'b1, 8'h9f, 8'h9e}; // CH=6 OP=3
cfg[3623] = { 1'b0, 8'h82, 8'h17}; // CH=2 OP=0
cfg[3624] = { 1'b1, 8'hfa, 8'hb1}; // CH=5 OP=2
cfg[3625] = { 1'b0, 8'hfc, 8'h45}; // CH=0 OP=3
cfg[3626] = { 1'b0, 8'h42, 8'h4e}; // CH=2 OP=0
cfg[3627] = { 1'b0, 8'hec, 8'h36}; // CH=0 OP=3
cfg[3628] = { 1'b1, 8'had, 8'h3e}; // CH=4 OP=3
cfg[3629] = { 1'b0, 8'h9c, 8'h88}; // CH=0 OP=3
cfg[3630] = { 1'b0, 8'h32, 8'h8d}; // CH=2 OP=0
cfg[3631] = { 1'b0, 8'hb4, 8'hde}; // CH=0 OP=1
cfg[3632] = { 1'b0, 8'hed, 8'h7e}; // CH=1 OP=3
cfg[3633] = { 1'b1, 8'h4b, 8'hfb}; // CH=6 OP=2
cfg[3634] = { 1'b0, 8'h87, 8'hf7}; // CH=3 OP=1
cfg[3635] = { 1'b0, 8'h77, 8'h3a}; // CH=3 OP=1
cfg[3636] = { 1'b0, 8'hd5, 8'h26}; // CH=1 OP=1
cfg[3637] = { 1'b0, 8'hef, 8'hd4}; // CH=3 OP=3
cfg[3638] = { 1'b1, 8'hfa, 8'h70}; // CH=5 OP=2
cfg[3639] = { 1'b1, 8'hf3, 8'h15}; // CH=6 OP=0
cfg[3640] = { 1'b1, 8'h71, 8'h1c}; // CH=4 OP=0
cfg[3641] = { 1'b1, 8'h72, 8'h48}; // CH=5 OP=0
cfg[3642] = { 1'b0, 8'h6d, 8'h25}; // CH=1 OP=3
cfg[3643] = { 1'b0, 8'h64, 8'h48}; // CH=0 OP=1
cfg[3644] = { 1'b1, 8'h9e, 8'hb8}; // CH=5 OP=3
cfg[3645] = { 1'b1, 8'hc5, 8'h5f}; // CH=4 OP=1
cfg[3646] = { 1'b0, 8'h99, 8'h43}; // CH=1 OP=2
cfg[3647] = { 1'b1, 8'hed, 8'hb0}; // CH=4 OP=3
cfg[3648] = { 1'b1, 8'hd8, 8'h9a}; // CH=3 OP=2
cfg[3649] = { 1'b0, 8'hb9, 8'hf6}; // CH=1 OP=2
cfg[3650] = { 1'b1, 8'ha6, 8'h67}; // CH=5 OP=1
cfg[3651] = { 1'b1, 8'h80, 8'hd9}; // CH=3 OP=0
cfg[3652] = { 1'b1, 8'ha6, 8'h46}; // CH=5 OP=1
cfg[3653] = { 1'b1, 8'h54, 8'hab}; // CH=3 OP=1
cfg[3654] = { 1'b1, 8'h79, 8'h49}; // CH=4 OP=2
cfg[3655] = { 1'b0, 8'h73, 8'he}; // CH=3 OP=0
cfg[3656] = { 1'b0, 8'h5c, 8'ha7}; // CH=0 OP=3
cfg[3657] = { 1'b0, 8'h4a, 8'hb0}; // CH=2 OP=2
cfg[3658] = { 1'b1, 8'h4c, 8'h4b}; // CH=3 OP=3
cfg[3659] = { 1'b1, 8'h42, 8'hed}; // CH=5 OP=0
cfg[3660] = { 1'b0, 8'haa, 8'hac}; // CH=2 OP=2
cfg[3661] = { 1'b0, 8'h83, 8'hb4}; // CH=3 OP=0
cfg[3662] = { 1'b1, 8'hca, 8'he1}; // CH=5 OP=2
cfg[3663] = { 1'b1, 8'h75, 8'h56}; // CH=4 OP=1
cfg[3664] = { 1'b1, 8'hbe, 8'h83}; // CH=5 OP=3
cfg[3665] = { 1'b0, 8'hcd, 8'h10}; // CH=1 OP=3
cfg[3666] = { 1'b1, 8'h74, 8'he0}; // CH=3 OP=1
cfg[3667] = { 1'b0, 8'h70, 8'h60}; // CH=0 OP=0
cfg[3668] = { 1'b0, 8'hbc, 8'h70}; // CH=0 OP=3
cfg[3669] = { 1'b1, 8'hff, 8'h5d}; // CH=6 OP=3
cfg[3670] = { 1'b0, 8'ha9, 8'ha}; // CH=1 OP=2
cfg[3671] = { 1'b0, 8'h91, 8'hbe}; // CH=1 OP=0
cfg[3672] = { 1'b1, 8'hf5, 8'hf6}; // CH=4 OP=1
cfg[3673] = { 1'b1, 8'h78, 8'hf8}; // CH=3 OP=2
cfg[3674] = { 1'b0, 8'h88, 8'h4f}; // CH=0 OP=2
cfg[3675] = { 1'b1, 8'h68, 8'h18}; // CH=3 OP=2
cfg[3676] = { 1'b1, 8'hc9, 8'h3e}; // CH=4 OP=2
cfg[3677] = { 1'b0, 8'h55, 8'hae}; // CH=1 OP=1
cfg[3678] = { 1'b0, 8'he4, 8'h6b}; // CH=0 OP=1
cfg[3679] = { 1'b0, 8'h30, 8'h6a}; // CH=0 OP=0
cfg[3680] = { 1'b0, 8'hdf, 8'h13}; // CH=3 OP=3
cfg[3681] = { 1'b0, 8'h70, 8'h3f}; // CH=0 OP=0
cfg[3682] = { 1'b1, 8'h8b, 8'h36}; // CH=6 OP=2
cfg[3683] = { 1'b0, 8'h84, 8'ha1}; // CH=0 OP=1
cfg[3684] = { 1'b0, 8'hd3, 8'hcb}; // CH=3 OP=0
cfg[3685] = { 1'b1, 8'heb, 8'hc2}; // CH=6 OP=2
cfg[3686] = { 1'b1, 8'hec, 8'h2e}; // CH=3 OP=3
cfg[3687] = { 1'b0, 8'h41, 8'hd8}; // CH=1 OP=0
cfg[3688] = { 1'b1, 8'had, 8'h43}; // CH=4 OP=3
cfg[3689] = { 1'b0, 8'hc0, 8'h85}; // CH=0 OP=0
cfg[3690] = { 1'b1, 8'ha6, 8'hab}; // CH=5 OP=1
cfg[3691] = { 1'b0, 8'h31, 8'h36}; // CH=1 OP=0
cfg[3692] = { 1'b0, 8'hb5, 8'hd7}; // CH=1 OP=1
cfg[3693] = { 1'b0, 8'h88, 8'ha3}; // CH=0 OP=2
cfg[3694] = { 1'b1, 8'h74, 8'h65}; // CH=3 OP=1
cfg[3695] = { 1'b1, 8'h9e, 8'h93}; // CH=5 OP=3
cfg[3696] = { 1'b1, 8'h76, 8'h52}; // CH=5 OP=1
cfg[3697] = { 1'b1, 8'hba, 8'h11}; // CH=5 OP=2
cfg[3698] = { 1'b1, 8'h67, 8'h2e}; // CH=6 OP=1
cfg[3699] = { 1'b1, 8'h5e, 8'hb3}; // CH=5 OP=3
cfg[3700] = { 1'b0, 8'hce, 8'hc1}; // CH=2 OP=3
cfg[3701] = { 1'b0, 8'hf8, 8'hf2}; // CH=0 OP=2
cfg[3702] = { 1'b1, 8'h54, 8'ha8}; // CH=3 OP=1
cfg[3703] = { 1'b0, 8'h6c, 8'h30}; // CH=0 OP=3
cfg[3704] = { 1'b0, 8'ha7, 8'ha4}; // CH=3 OP=1
cfg[3705] = { 1'b1, 8'hce, 8'h42}; // CH=5 OP=3
cfg[3706] = { 1'b1, 8'h37, 8'hb9}; // CH=6 OP=1
cfg[3707] = { 1'b0, 8'hc6, 8'h73}; // CH=2 OP=1
cfg[3708] = { 1'b0, 8'hac, 8'hda}; // CH=0 OP=3
cfg[3709] = { 1'b1, 8'hc7, 8'h2}; // CH=6 OP=1
cfg[3710] = { 1'b1, 8'h88, 8'h2a}; // CH=3 OP=2
cfg[3711] = { 1'b1, 8'h7a, 8'h88}; // CH=5 OP=2
cfg[3712] = { 1'b1, 8'h8e, 8'hbe}; // CH=5 OP=3
cfg[3713] = { 1'b0, 8'hfa, 8'h53}; // CH=2 OP=2
cfg[3714] = { 1'b0, 8'ha1, 8'hf7}; // CH=1 OP=0
cfg[3715] = { 1'b0, 8'h6f, 8'h3a}; // CH=3 OP=3
cfg[3716] = { 1'b1, 8'ha7, 8'hf3}; // CH=6 OP=1
cfg[3717] = { 1'b0, 8'h6d, 8'h66}; // CH=1 OP=3
cfg[3718] = { 1'b0, 8'h76, 8'h40}; // CH=2 OP=1
cfg[3719] = { 1'b1, 8'he9, 8'he0}; // CH=4 OP=2
cfg[3720] = { 1'b1, 8'hf6, 8'h68}; // CH=5 OP=1
cfg[3721] = { 1'b1, 8'hb4, 8'h64}; // CH=3 OP=1
cfg[3722] = { 1'b1, 8'h4a, 8'hf2}; // CH=5 OP=2
cfg[3723] = { 1'b0, 8'h50, 8'hec}; // CH=0 OP=0
cfg[3724] = { 1'b1, 8'h8a, 8'hc5}; // CH=5 OP=2
cfg[3725] = { 1'b1, 8'h7d, 8'h8e}; // CH=4 OP=3
cfg[3726] = { 1'b0, 8'he3, 8'h8c}; // CH=3 OP=0
cfg[3727] = { 1'b1, 8'h63, 8'hed}; // CH=6 OP=0
cfg[3728] = { 1'b0, 8'h4c, 8'hb}; // CH=0 OP=3
cfg[3729] = { 1'b0, 8'h77, 8'h74}; // CH=3 OP=1
cfg[3730] = { 1'b0, 8'hdc, 8'h57}; // CH=0 OP=3
cfg[3731] = { 1'b0, 8'hce, 8'h5c}; // CH=2 OP=3
cfg[3732] = { 1'b0, 8'hbb, 8'hb5}; // CH=3 OP=2
cfg[3733] = { 1'b1, 8'h48, 8'h5}; // CH=3 OP=2
cfg[3734] = { 1'b0, 8'h45, 8'h8f}; // CH=1 OP=1
cfg[3735] = { 1'b1, 8'he9, 8'hc}; // CH=4 OP=2
cfg[3736] = { 1'b1, 8'hfb, 8'hef}; // CH=6 OP=2
cfg[3737] = { 1'b0, 8'h79, 8'h12}; // CH=1 OP=2
cfg[3738] = { 1'b1, 8'h4d, 8'h64}; // CH=4 OP=3
cfg[3739] = { 1'b1, 8'hfc, 8'hdb}; // CH=3 OP=3
cfg[3740] = { 1'b1, 8'h59, 8'h95}; // CH=4 OP=2
cfg[3741] = { 1'b0, 8'h41, 8'h5d}; // CH=1 OP=0
cfg[3742] = { 1'b1, 8'h89, 8'h13}; // CH=4 OP=2
cfg[3743] = { 1'b1, 8'hcf, 8'ha2}; // CH=6 OP=3
cfg[3744] = { 1'b0, 8'hb8, 8'hae}; // CH=0 OP=2
cfg[3745] = { 1'b0, 8'hb3, 8'h9d}; // CH=3 OP=0
cfg[3746] = { 1'b0, 8'hd9, 8'haf}; // CH=1 OP=2
cfg[3747] = { 1'b0, 8'h75, 8'h28}; // CH=1 OP=1
cfg[3748] = { 1'b0, 8'h8c, 8'hff}; // CH=0 OP=3
cfg[3749] = { 1'b1, 8'h3d, 8'hb7}; // CH=4 OP=3
cfg[3750] = { 1'b1, 8'h7e, 8'h14}; // CH=5 OP=3
cfg[3751] = { 1'b0, 8'hb5, 8'h27}; // CH=1 OP=1
cfg[3752] = { 1'b1, 8'he2, 8'hd6}; // CH=5 OP=0
cfg[3753] = { 1'b1, 8'hd6, 8'h8f}; // CH=5 OP=1
cfg[3754] = { 1'b0, 8'h7e, 8'h42}; // CH=2 OP=3
cfg[3755] = { 1'b1, 8'h3e, 8'h1c}; // CH=5 OP=3
cfg[3756] = { 1'b0, 8'h62, 8'h27}; // CH=2 OP=0
cfg[3757] = { 1'b1, 8'h62, 8'hd7}; // CH=5 OP=0
cfg[3758] = { 1'b0, 8'h8a, 8'h84}; // CH=2 OP=2
cfg[3759] = { 1'b0, 8'h9e, 8'h8e}; // CH=2 OP=3
cfg[3760] = { 1'b0, 8'hc5, 8'h52}; // CH=1 OP=1
cfg[3761] = { 1'b1, 8'h8e, 8'h8}; // CH=5 OP=3
cfg[3762] = { 1'b0, 8'h41, 8'hea}; // CH=1 OP=0
cfg[3763] = { 1'b0, 8'h83, 8'h19}; // CH=3 OP=0
cfg[3764] = { 1'b0, 8'h9f, 8'hdd}; // CH=3 OP=3
cfg[3765] = { 1'b1, 8'hc6, 8'hc9}; // CH=5 OP=1
cfg[3766] = { 1'b1, 8'h9e, 8'h2a}; // CH=5 OP=3
cfg[3767] = { 1'b1, 8'h5a, 8'h18}; // CH=5 OP=2
cfg[3768] = { 1'b0, 8'hb0, 8'had}; // CH=0 OP=0
cfg[3769] = { 1'b0, 8'h84, 8'h4b}; // CH=0 OP=1
cfg[3770] = { 1'b1, 8'h60, 8'h11}; // CH=3 OP=0
cfg[3771] = { 1'b1, 8'hfb, 8'h9f}; // CH=6 OP=2
cfg[3772] = { 1'b1, 8'hbb, 8'h53}; // CH=6 OP=2
cfg[3773] = { 1'b0, 8'hf9, 8'hd6}; // CH=1 OP=2
cfg[3774] = { 1'b1, 8'h76, 8'h76}; // CH=5 OP=1
cfg[3775] = { 1'b0, 8'h56, 8'h3c}; // CH=2 OP=1
cfg[3776] = { 1'b1, 8'h97, 8'hda}; // CH=6 OP=1
cfg[3777] = { 1'b1, 8'hf2, 8'hfd}; // CH=5 OP=0
cfg[3778] = { 1'b1, 8'ha2, 8'haa}; // CH=5 OP=0
cfg[3779] = { 1'b0, 8'h8f, 8'hf5}; // CH=3 OP=3
cfg[3780] = { 1'b0, 8'ha0, 8'h87}; // CH=0 OP=0
cfg[3781] = { 1'b0, 8'h9b, 8'h99}; // CH=3 OP=2
cfg[3782] = { 1'b1, 8'h56, 8'hec}; // CH=5 OP=1
cfg[3783] = { 1'b1, 8'h4f, 8'hc2}; // CH=6 OP=3
cfg[3784] = { 1'b1, 8'hc6, 8'h38}; // CH=5 OP=1
cfg[3785] = { 1'b1, 8'h98, 8'h75}; // CH=3 OP=2
cfg[3786] = { 1'b1, 8'h40, 8'hb3}; // CH=3 OP=0
cfg[3787] = { 1'b0, 8'hf6, 8'ha5}; // CH=2 OP=1
cfg[3788] = { 1'b0, 8'hec, 8'h95}; // CH=0 OP=3
cfg[3789] = { 1'b1, 8'hf2, 8'h24}; // CH=5 OP=0
cfg[3790] = { 1'b0, 8'h98, 8'hc4}; // CH=0 OP=2
cfg[3791] = { 1'b1, 8'he3, 8'h5f}; // CH=6 OP=0
cfg[3792] = { 1'b1, 8'hed, 8'hb5}; // CH=4 OP=3
cfg[3793] = { 1'b1, 8'h92, 8'h5}; // CH=5 OP=0
cfg[3794] = { 1'b0, 8'h9b, 8'hcb}; // CH=3 OP=2
cfg[3795] = { 1'b1, 8'h34, 8'he7}; // CH=3 OP=1
cfg[3796] = { 1'b0, 8'h74, 8'h9a}; // CH=0 OP=1
cfg[3797] = { 1'b1, 8'h83, 8'h40}; // CH=6 OP=0
cfg[3798] = { 1'b1, 8'h69, 8'h88}; // CH=4 OP=2
cfg[3799] = { 1'b1, 8'h5c, 8'h3d}; // CH=3 OP=3
cfg[3800] = { 1'b1, 8'hf4, 8'h2}; // CH=3 OP=1
cfg[3801] = { 1'b0, 8'hd8, 8'h61}; // CH=0 OP=2
cfg[3802] = { 1'b1, 8'hc5, 8'h17}; // CH=4 OP=1
cfg[3803] = { 1'b0, 8'h57, 8'h1c}; // CH=3 OP=1
cfg[3804] = { 1'b0, 8'hf2, 8'he7}; // CH=2 OP=0
cfg[3805] = { 1'b1, 8'hd0, 8'hce}; // CH=3 OP=0
cfg[3806] = { 1'b0, 8'h57, 8'h9a}; // CH=3 OP=1
cfg[3807] = { 1'b0, 8'hd4, 8'h1e}; // CH=0 OP=1
cfg[3808] = { 1'b0, 8'h3e, 8'h37}; // CH=2 OP=3
cfg[3809] = { 1'b1, 8'h9a, 8'h74}; // CH=5 OP=2
cfg[3810] = { 1'b0, 8'h8e, 8'h76}; // CH=2 OP=3
cfg[3811] = { 1'b0, 8'h66, 8'hd8}; // CH=2 OP=1
cfg[3812] = { 1'b1, 8'hbc, 8'hef}; // CH=3 OP=3
cfg[3813] = { 1'b1, 8'h66, 8'h82}; // CH=5 OP=1
cfg[3814] = { 1'b0, 8'hfc, 8'h75}; // CH=0 OP=3
cfg[3815] = { 1'b0, 8'hcc, 8'h9b}; // CH=0 OP=3
cfg[3816] = { 1'b0, 8'hd1, 8'h36}; // CH=1 OP=0
cfg[3817] = { 1'b0, 8'h8b, 8'hf7}; // CH=3 OP=2
cfg[3818] = { 1'b1, 8'hff, 8'h29}; // CH=6 OP=3
cfg[3819] = { 1'b1, 8'h76, 8'h3d}; // CH=5 OP=1
cfg[3820] = { 1'b0, 8'h4e, 8'hce}; // CH=2 OP=3
cfg[3821] = { 1'b0, 8'h3d, 8'h55}; // CH=1 OP=3
cfg[3822] = { 1'b0, 8'h48, 8'h11}; // CH=0 OP=2
cfg[3823] = { 1'b0, 8'h3a, 8'h78}; // CH=2 OP=2
cfg[3824] = { 1'b1, 8'hfa, 8'h74}; // CH=5 OP=2
cfg[3825] = { 1'b1, 8'hb9, 8'h40}; // CH=4 OP=2
cfg[3826] = { 1'b1, 8'h5a, 8'hf3}; // CH=5 OP=2
cfg[3827] = { 1'b1, 8'h90, 8'h98}; // CH=3 OP=0
cfg[3828] = { 1'b0, 8'h5f, 8'h97}; // CH=3 OP=3
cfg[3829] = { 1'b1, 8'hbd, 8'hd}; // CH=4 OP=3
cfg[3830] = { 1'b1, 8'h82, 8'h5b}; // CH=5 OP=0
cfg[3831] = { 1'b1, 8'h72, 8'h98}; // CH=5 OP=0
cfg[3832] = { 1'b0, 8'he4, 8'he0}; // CH=0 OP=1
cfg[3833] = { 1'b0, 8'hcc, 8'h1a}; // CH=0 OP=3
cfg[3834] = { 1'b0, 8'h4f, 8'h14}; // CH=3 OP=3
cfg[3835] = { 1'b0, 8'h7a, 8'h37}; // CH=2 OP=2
cfg[3836] = { 1'b1, 8'h3d, 8'had}; // CH=4 OP=3
cfg[3837] = { 1'b0, 8'h99, 8'h69}; // CH=1 OP=2
cfg[3838] = { 1'b0, 8'hc2, 8'h27}; // CH=2 OP=0
cfg[3839] = { 1'b1, 8'h41, 8'ha9}; // CH=4 OP=0
cfg[3840] = { 1'b0, 8'hd2, 8'h1b}; // CH=2 OP=0
cfg[3841] = { 1'b0, 8'hda, 8'hff}; // CH=2 OP=2
cfg[3842] = { 1'b1, 8'h57, 8'hcb}; // CH=6 OP=1
cfg[3843] = { 1'b1, 8'h8c, 8'h1a}; // CH=3 OP=3
cfg[3844] = { 1'b0, 8'hb7, 8'h33}; // CH=3 OP=1
cfg[3845] = { 1'b1, 8'hd6, 8'had}; // CH=5 OP=1
cfg[3846] = { 1'b0, 8'had, 8'hb7}; // CH=1 OP=3
cfg[3847] = { 1'b1, 8'h6f, 8'h47}; // CH=6 OP=3
cfg[3848] = { 1'b0, 8'hb1, 8'hf0}; // CH=1 OP=0
cfg[3849] = { 1'b0, 8'h83, 8'hb}; // CH=3 OP=0
cfg[3850] = { 1'b1, 8'h5d, 8'hb}; // CH=4 OP=3
cfg[3851] = { 1'b0, 8'hb4, 8'hd6}; // CH=0 OP=1
cfg[3852] = { 1'b1, 8'hc8, 8'hf1}; // CH=3 OP=2
cfg[3853] = { 1'b0, 8'hfb, 8'h13}; // CH=3 OP=2
cfg[3854] = { 1'b1, 8'ha8, 8'h4b}; // CH=3 OP=2
cfg[3855] = { 1'b1, 8'h5f, 8'h2f}; // CH=6 OP=3
cfg[3856] = { 1'b1, 8'h7f, 8'h58}; // CH=6 OP=3
cfg[3857] = { 1'b0, 8'hc7, 8'hd3}; // CH=3 OP=1
cfg[3858] = { 1'b0, 8'hb7, 8'hfc}; // CH=3 OP=1
cfg[3859] = { 1'b1, 8'hc3, 8'h6a}; // CH=6 OP=0
cfg[3860] = { 1'b0, 8'hce, 8'hff}; // CH=2 OP=3
cfg[3861] = { 1'b1, 8'ha4, 8'hd5}; // CH=3 OP=1
cfg[3862] = { 1'b0, 8'h95, 8'h1}; // CH=1 OP=1
cfg[3863] = { 1'b0, 8'ha9, 8'hb9}; // CH=1 OP=2
cfg[3864] = { 1'b1, 8'hf4, 8'h28}; // CH=3 OP=1
cfg[3865] = { 1'b1, 8'h86, 8'h6d}; // CH=5 OP=1
cfg[3866] = { 1'b1, 8'hcd, 8'h7c}; // CH=4 OP=3
cfg[3867] = { 1'b1, 8'h43, 8'hcc}; // CH=6 OP=0
cfg[3868] = { 1'b1, 8'h6a, 8'h84}; // CH=5 OP=2
cfg[3869] = { 1'b0, 8'hb5, 8'h47}; // CH=1 OP=1
cfg[3870] = { 1'b1, 8'h8b, 8'h1c}; // CH=6 OP=2
cfg[3871] = { 1'b1, 8'h8c, 8'hd8}; // CH=3 OP=3
cfg[3872] = { 1'b1, 8'h45, 8'h5c}; // CH=4 OP=1
cfg[3873] = { 1'b0, 8'h6d, 8'hdb}; // CH=1 OP=3
cfg[3874] = { 1'b0, 8'hda, 8'h2}; // CH=2 OP=2
cfg[3875] = { 1'b1, 8'ha1, 8'h88}; // CH=4 OP=0
cfg[3876] = { 1'b1, 8'h6f, 8'h8d}; // CH=6 OP=3
cfg[3877] = { 1'b1, 8'hb2, 8'h5a}; // CH=5 OP=0
cfg[3878] = { 1'b0, 8'hdc, 8'hde}; // CH=0 OP=3
cfg[3879] = { 1'b1, 8'h92, 8'h31}; // CH=5 OP=0
cfg[3880] = { 1'b0, 8'hf3, 8'h4d}; // CH=3 OP=0
cfg[3881] = { 1'b1, 8'h42, 8'ha9}; // CH=5 OP=0
cfg[3882] = { 1'b1, 8'h3a, 8'hee}; // CH=5 OP=2
cfg[3883] = { 1'b0, 8'h5e, 8'h5b}; // CH=2 OP=3
cfg[3884] = { 1'b1, 8'he6, 8'h36}; // CH=5 OP=1
cfg[3885] = { 1'b1, 8'h74, 8'hc1}; // CH=3 OP=1
cfg[3886] = { 1'b0, 8'hce, 8'h9c}; // CH=2 OP=3
cfg[3887] = { 1'b0, 8'hac, 8'hc3}; // CH=0 OP=3
cfg[3888] = { 1'b1, 8'hd1, 8'h9f}; // CH=4 OP=0
cfg[3889] = { 1'b1, 8'h94, 8'h31}; // CH=3 OP=1
cfg[3890] = { 1'b0, 8'hba, 8'hfe}; // CH=2 OP=2
cfg[3891] = { 1'b1, 8'h3b, 8'h41}; // CH=6 OP=2
cfg[3892] = { 1'b1, 8'h98, 8'h7b}; // CH=3 OP=2
cfg[3893] = { 1'b0, 8'hf6, 8'ha2}; // CH=2 OP=1
cfg[3894] = { 1'b0, 8'hdd, 8'hd8}; // CH=1 OP=3
cfg[3895] = { 1'b1, 8'h51, 8'h99}; // CH=4 OP=0
cfg[3896] = { 1'b1, 8'h8b, 8'h36}; // CH=6 OP=2
cfg[3897] = { 1'b1, 8'ha1, 8'hcb}; // CH=4 OP=0
cfg[3898] = { 1'b0, 8'he8, 8'h9c}; // CH=0 OP=2
cfg[3899] = { 1'b0, 8'h7c, 8'ha7}; // CH=0 OP=3
cfg[3900] = { 1'b0, 8'h36, 8'ha5}; // CH=2 OP=1
cfg[3901] = { 1'b0, 8'h72, 8'he6}; // CH=2 OP=0
cfg[3902] = { 1'b1, 8'h36, 8'h62}; // CH=5 OP=1
cfg[3903] = { 1'b0, 8'hac, 8'h0}; // CH=0 OP=3
cfg[3904] = { 1'b0, 8'hf9, 8'hdd}; // CH=1 OP=2
cfg[3905] = { 1'b1, 8'h8c, 8'h2e}; // CH=3 OP=3
cfg[3906] = { 1'b1, 8'ha4, 8'h4d}; // CH=3 OP=1
cfg[3907] = { 1'b0, 8'h3d, 8'hb8}; // CH=1 OP=3
cfg[3908] = { 1'b0, 8'h5b, 8'ha0}; // CH=3 OP=2
cfg[3909] = { 1'b1, 8'h53, 8'h1f}; // CH=6 OP=0
cfg[3910] = { 1'b1, 8'hc5, 8'he7}; // CH=4 OP=1
cfg[3911] = { 1'b1, 8'hcf, 8'h49}; // CH=6 OP=3
cfg[3912] = { 1'b1, 8'hd0, 8'h4d}; // CH=3 OP=0
cfg[3913] = { 1'b1, 8'had, 8'h29}; // CH=4 OP=3
cfg[3914] = { 1'b0, 8'hdc, 8'h9f}; // CH=0 OP=3
cfg[3915] = { 1'b0, 8'ha3, 8'h4a}; // CH=3 OP=0
cfg[3916] = { 1'b1, 8'h5c, 8'h42}; // CH=3 OP=3
cfg[3917] = { 1'b0, 8'hfc, 8'hf6}; // CH=0 OP=3
cfg[3918] = { 1'b1, 8'h52, 8'h52}; // CH=5 OP=0
cfg[3919] = { 1'b1, 8'h82, 8'h6d}; // CH=5 OP=0
cfg[3920] = { 1'b0, 8'ha7, 8'h32}; // CH=3 OP=1
cfg[3921] = { 1'b0, 8'hd1, 8'h2}; // CH=1 OP=0
cfg[3922] = { 1'b0, 8'hfb, 8'h9}; // CH=3 OP=2
cfg[3923] = { 1'b1, 8'h9a, 8'h9}; // CH=5 OP=2
cfg[3924] = { 1'b1, 8'he4, 8'h95}; // CH=3 OP=1
cfg[3925] = { 1'b1, 8'hd3, 8'h38}; // CH=6 OP=0
cfg[3926] = { 1'b1, 8'hff, 8'h94}; // CH=6 OP=3
cfg[3927] = { 1'b1, 8'h32, 8'h91}; // CH=5 OP=0
cfg[3928] = { 1'b1, 8'h85, 8'haa}; // CH=4 OP=1
cfg[3929] = { 1'b0, 8'h9d, 8'h17}; // CH=1 OP=3
cfg[3930] = { 1'b0, 8'h4c, 8'hae}; // CH=0 OP=3
cfg[3931] = { 1'b0, 8'hb9, 8'hf2}; // CH=1 OP=2
cfg[3932] = { 1'b1, 8'hc2, 8'h9d}; // CH=5 OP=0
cfg[3933] = { 1'b1, 8'h57, 8'hf9}; // CH=6 OP=1
cfg[3934] = { 1'b0, 8'h8f, 8'h7e}; // CH=3 OP=3
cfg[3935] = { 1'b1, 8'h3f, 8'h45}; // CH=6 OP=3
cfg[3936] = { 1'b0, 8'h71, 8'hb5}; // CH=1 OP=0
cfg[3937] = { 1'b0, 8'hf6, 8'h5f}; // CH=2 OP=1
cfg[3938] = { 1'b0, 8'hfd, 8'h77}; // CH=1 OP=3
cfg[3939] = { 1'b1, 8'hab, 8'hc1}; // CH=6 OP=2
cfg[3940] = { 1'b0, 8'h5b, 8'hd}; // CH=3 OP=2
cfg[3941] = { 1'b1, 8'hc8, 8'h2b}; // CH=3 OP=2
cfg[3942] = { 1'b0, 8'hc1, 8'h9a}; // CH=1 OP=0
cfg[3943] = { 1'b1, 8'h3f, 8'h6}; // CH=6 OP=3
cfg[3944] = { 1'b1, 8'h84, 8'h45}; // CH=3 OP=1
cfg[3945] = { 1'b1, 8'h87, 8'h84}; // CH=6 OP=1
cfg[3946] = { 1'b0, 8'h99, 8'hf6}; // CH=1 OP=2
cfg[3947] = { 1'b1, 8'h6c, 8'hec}; // CH=3 OP=3
cfg[3948] = { 1'b0, 8'h95, 8'h1f}; // CH=1 OP=1
cfg[3949] = { 1'b1, 8'hf1, 8'h3a}; // CH=4 OP=0
cfg[3950] = { 1'b0, 8'h89, 8'h65}; // CH=1 OP=2
cfg[3951] = { 1'b0, 8'hef, 8'hdc}; // CH=3 OP=3
cfg[3952] = { 1'b1, 8'hc6, 8'h29}; // CH=5 OP=1
cfg[3953] = { 1'b0, 8'ha7, 8'hb3}; // CH=3 OP=1
cfg[3954] = { 1'b1, 8'h3d, 8'h3a}; // CH=4 OP=3
cfg[3955] = { 1'b1, 8'h33, 8'hd3}; // CH=6 OP=0
cfg[3956] = { 1'b1, 8'h9f, 8'he1}; // CH=6 OP=3
cfg[3957] = { 1'b1, 8'hcd, 8'h0}; // CH=4 OP=3
cfg[3958] = { 1'b1, 8'h46, 8'h51}; // CH=5 OP=1
cfg[3959] = { 1'b0, 8'h4b, 8'h6d}; // CH=3 OP=2
cfg[3960] = { 1'b1, 8'h74, 8'h9b}; // CH=3 OP=1
cfg[3961] = { 1'b0, 8'h9d, 8'h31}; // CH=1 OP=3
cfg[3962] = { 1'b1, 8'h6d, 8'hf7}; // CH=4 OP=3
cfg[3963] = { 1'b1, 8'ha7, 8'hfe}; // CH=6 OP=1
cfg[3964] = { 1'b0, 8'h7b, 8'he7}; // CH=3 OP=2
cfg[3965] = { 1'b1, 8'h5c, 8'hbd}; // CH=3 OP=3
cfg[3966] = { 1'b1, 8'h5c, 8'h7c}; // CH=3 OP=3
cfg[3967] = { 1'b0, 8'had, 8'hd1}; // CH=1 OP=3
cfg[3968] = { 1'b1, 8'h75, 8'h17}; // CH=4 OP=1
cfg[3969] = { 1'b0, 8'hc6, 8'h63}; // CH=2 OP=1
cfg[3970] = { 1'b1, 8'h3a, 8'h8a}; // CH=5 OP=2
cfg[3971] = { 1'b0, 8'hd7, 8'hbb}; // CH=3 OP=1
cfg[3972] = { 1'b1, 8'he3, 8'hb3}; // CH=6 OP=0
cfg[3973] = { 1'b0, 8'he1, 8'h52}; // CH=1 OP=0
cfg[3974] = { 1'b0, 8'hc9, 8'h2e}; // CH=1 OP=2
cfg[3975] = { 1'b1, 8'h86, 8'h3e}; // CH=5 OP=1
cfg[3976] = { 1'b1, 8'h69, 8'hed}; // CH=4 OP=2
cfg[3977] = { 1'b0, 8'hec, 8'hc4}; // CH=0 OP=3
cfg[3978] = { 1'b1, 8'hdd, 8'h3a}; // CH=4 OP=3
cfg[3979] = { 1'b0, 8'h68, 8'h0}; // CH=0 OP=2
cfg[3980] = { 1'b1, 8'h7e, 8'h3b}; // CH=5 OP=3
cfg[3981] = { 1'b0, 8'h4e, 8'h12}; // CH=2 OP=3
cfg[3982] = { 1'b1, 8'h8a, 8'hf5}; // CH=5 OP=2
cfg[3983] = { 1'b1, 8'h6e, 8'hd7}; // CH=5 OP=3
cfg[3984] = { 1'b0, 8'hcd, 8'ha0}; // CH=1 OP=3
cfg[3985] = { 1'b0, 8'h88, 8'h26}; // CH=0 OP=2
cfg[3986] = { 1'b1, 8'h9f, 8'h28}; // CH=6 OP=3
cfg[3987] = { 1'b0, 8'h64, 8'hfc}; // CH=0 OP=1
cfg[3988] = { 1'b0, 8'h9e, 8'he8}; // CH=2 OP=3
cfg[3989] = { 1'b1, 8'h9e, 8'h36}; // CH=5 OP=3
cfg[3990] = { 1'b0, 8'hd9, 8'hf}; // CH=1 OP=2
cfg[3991] = { 1'b0, 8'hec, 8'ha4}; // CH=0 OP=3
cfg[3992] = { 1'b0, 8'he1, 8'heb}; // CH=1 OP=0
cfg[3993] = { 1'b1, 8'hb8, 8'h85}; // CH=3 OP=2
cfg[3994] = { 1'b1, 8'h58, 8'h4d}; // CH=3 OP=2
cfg[3995] = { 1'b1, 8'h7e, 8'h53}; // CH=5 OP=3
cfg[3996] = { 1'b1, 8'ha7, 8'h46}; // CH=6 OP=1
cfg[3997] = { 1'b1, 8'ha3, 8'ha2}; // CH=6 OP=0
cfg[3998] = { 1'b1, 8'h8b, 8'hea}; // CH=6 OP=2
cfg[3999] = { 1'b1, 8'hc2, 8'h10}; // CH=5 OP=0
cfg[4000] = { 1'b1, 8'hd1, 8'h9e}; // CH=4 OP=0
cfg[4001] = { 1'b1, 8'h75, 8'haa}; // CH=4 OP=1
cfg[4002] = { 1'b1, 8'h61, 8'h5}; // CH=4 OP=0
cfg[4003] = { 1'b0, 8'he6, 8'hea}; // CH=2 OP=1
cfg[4004] = { 1'b1, 8'h33, 8'h3d}; // CH=6 OP=0
cfg[4005] = { 1'b1, 8'h86, 8'h5e}; // CH=5 OP=1
cfg[4006] = { 1'b0, 8'hcc, 8'h8}; // CH=0 OP=3
cfg[4007] = { 1'b1, 8'h6e, 8'h51}; // CH=5 OP=3
cfg[4008] = { 1'b0, 8'h58, 8'hfe}; // CH=0 OP=2
cfg[4009] = { 1'b0, 8'h68, 8'h49}; // CH=0 OP=2
cfg[4010] = { 1'b0, 8'h89, 8'h32}; // CH=1 OP=2
cfg[4011] = { 1'b1, 8'hff, 8'hb1}; // CH=6 OP=3
cfg[4012] = { 1'b0, 8'h60, 8'hb6}; // CH=0 OP=0
cfg[4013] = { 1'b1, 8'h46, 8'ha0}; // CH=5 OP=1
cfg[4014] = { 1'b0, 8'h79, 8'hdd}; // CH=1 OP=2
cfg[4015] = { 1'b1, 8'hff, 8'h3c}; // CH=6 OP=3
cfg[4016] = { 1'b1, 8'hcb, 8'h44}; // CH=6 OP=2
cfg[4017] = { 1'b0, 8'h39, 8'h95}; // CH=1 OP=2
cfg[4018] = { 1'b1, 8'h91, 8'h93}; // CH=4 OP=0
cfg[4019] = { 1'b1, 8'hfa, 8'hdc}; // CH=5 OP=2
cfg[4020] = { 1'b1, 8'ha8, 8'he}; // CH=3 OP=2
cfg[4021] = { 1'b0, 8'ha7, 8'hb1}; // CH=3 OP=1
cfg[4022] = { 1'b0, 8'hdd, 8'h67}; // CH=1 OP=3
cfg[4023] = { 1'b1, 8'h5b, 8'h4d}; // CH=6 OP=2
cfg[4024] = { 1'b1, 8'h7b, 8'hc6}; // CH=6 OP=2
cfg[4025] = { 1'b1, 8'hba, 8'hc5}; // CH=5 OP=2
cfg[4026] = { 1'b1, 8'hc1, 8'h90}; // CH=4 OP=0
cfg[4027] = { 1'b0, 8'h32, 8'hc9}; // CH=2 OP=0
cfg[4028] = { 1'b1, 8'h99, 8'h5b}; // CH=4 OP=2
cfg[4029] = { 1'b1, 8'hb8, 8'h55}; // CH=3 OP=2
cfg[4030] = { 1'b1, 8'h60, 8'h55}; // CH=3 OP=0
cfg[4031] = { 1'b1, 8'h6e, 8'h7}; // CH=5 OP=3
cfg[4032] = { 1'b1, 8'h76, 8'h1}; // CH=5 OP=1
cfg[4033] = { 1'b1, 8'h5b, 8'h5d}; // CH=6 OP=2
cfg[4034] = { 1'b1, 8'h7c, 8'hd8}; // CH=3 OP=3
cfg[4035] = { 1'b1, 8'he1, 8'h92}; // CH=4 OP=0
cfg[4036] = { 1'b1, 8'hdb, 8'h53}; // CH=6 OP=2
cfg[4037] = { 1'b1, 8'h68, 8'h85}; // CH=3 OP=2
cfg[4038] = { 1'b0, 8'hd1, 8'h1e}; // CH=1 OP=0
cfg[4039] = { 1'b1, 8'h48, 8'hd6}; // CH=3 OP=2
cfg[4040] = { 1'b0, 8'hc4, 8'h37}; // CH=0 OP=1
cfg[4041] = { 1'b1, 8'he8, 8'h3f}; // CH=3 OP=2
cfg[4042] = { 1'b0, 8'he9, 8'h4e}; // CH=1 OP=2
cfg[4043] = { 1'b0, 8'h46, 8'hab}; // CH=2 OP=1
cfg[4044] = { 1'b1, 8'hb8, 8'hcf}; // CH=3 OP=2
cfg[4045] = { 1'b1, 8'h31, 8'hec}; // CH=4 OP=0
cfg[4046] = { 1'b0, 8'h74, 8'hc7}; // CH=0 OP=1
cfg[4047] = { 1'b0, 8'ha8, 8'h2f}; // CH=0 OP=2
cfg[4048] = { 1'b0, 8'h7f, 8'h5}; // CH=3 OP=3
cfg[4049] = { 1'b0, 8'hb6, 8'h4e}; // CH=2 OP=1
cfg[4050] = { 1'b0, 8'hf5, 8'h9d}; // CH=1 OP=1
cfg[4051] = { 1'b0, 8'h43, 8'h5b}; // CH=3 OP=0
cfg[4052] = { 1'b0, 8'hef, 8'h8f}; // CH=3 OP=3
cfg[4053] = { 1'b0, 8'hbe, 8'h1e}; // CH=2 OP=3
cfg[4054] = { 1'b1, 8'h76, 8'h29}; // CH=5 OP=1
cfg[4055] = { 1'b0, 8'ha7, 8'h15}; // CH=3 OP=1
cfg[4056] = { 1'b0, 8'h82, 8'hdc}; // CH=2 OP=0
cfg[4057] = { 1'b1, 8'h34, 8'h2e}; // CH=3 OP=1
cfg[4058] = { 1'b0, 8'h82, 8'h54}; // CH=2 OP=0
cfg[4059] = { 1'b0, 8'h55, 8'h60}; // CH=1 OP=1
cfg[4060] = { 1'b1, 8'h98, 8'h7b}; // CH=3 OP=2
cfg[4061] = { 1'b1, 8'h87, 8'ha}; // CH=6 OP=1
cfg[4062] = { 1'b1, 8'h45, 8'h29}; // CH=4 OP=1
cfg[4063] = { 1'b0, 8'hbb, 8'h52}; // CH=3 OP=2
cfg[4064] = { 1'b0, 8'h63, 8'h68}; // CH=3 OP=0
cfg[4065] = { 1'b1, 8'h7f, 8'h44}; // CH=6 OP=3
cfg[4066] = { 1'b1, 8'had, 8'h50}; // CH=4 OP=3
cfg[4067] = { 1'b0, 8'he1, 8'h5b}; // CH=1 OP=0
cfg[4068] = { 1'b0, 8'h63, 8'haf}; // CH=3 OP=0
cfg[4069] = { 1'b0, 8'h83, 8'h10}; // CH=3 OP=0
cfg[4070] = { 1'b1, 8'hfe, 8'h65}; // CH=5 OP=3
cfg[4071] = { 1'b0, 8'hb3, 8'h98}; // CH=3 OP=0
cfg[4072] = { 1'b1, 8'hf9, 8'h31}; // CH=4 OP=2
cfg[4073] = { 1'b0, 8'hb4, 8'h84}; // CH=0 OP=1
cfg[4074] = { 1'b0, 8'h9f, 8'hec}; // CH=3 OP=3
cfg[4075] = { 1'b0, 8'ha9, 8'h96}; // CH=1 OP=2
cfg[4076] = { 1'b0, 8'hdd, 8'h44}; // CH=1 OP=3
cfg[4077] = { 1'b0, 8'hbc, 8'h25}; // CH=0 OP=3
cfg[4078] = { 1'b1, 8'hfa, 8'h89}; // CH=5 OP=2
cfg[4079] = { 1'b1, 8'h8e, 8'hc}; // CH=5 OP=3
cfg[4080] = { 1'b0, 8'hba, 8'ha}; // CH=2 OP=2
cfg[4081] = { 1'b0, 8'h6d, 8'h12}; // CH=1 OP=3
cfg[4082] = { 1'b0, 8'h66, 8'h44}; // CH=2 OP=1
cfg[4083] = { 1'b0, 8'hb4, 8'hc8}; // CH=0 OP=1
cfg[4084] = { 1'b0, 8'he4, 8'hca}; // CH=0 OP=1
cfg[4085] = { 1'b1, 8'h65, 8'h73}; // CH=4 OP=1
cfg[4086] = { 1'b1, 8'h41, 8'h50}; // CH=4 OP=0
cfg[4087] = { 1'b0, 8'hcc, 8'hc}; // CH=0 OP=3
cfg[4088] = { 1'b1, 8'h68, 8'h7}; // CH=3 OP=2
cfg[4089] = { 1'b1, 8'h68, 8'h95}; // CH=3 OP=2
cfg[4090] = { 1'b1, 8'he4, 8'h4f}; // CH=3 OP=1
cfg[4091] = { 1'b0, 8'h9b, 8'h89}; // CH=3 OP=2
cfg[4092] = { 1'b0, 8'hc5, 8'h3e}; // CH=1 OP=1
cfg[4093] = { 1'b0, 8'h8f, 8'h70}; // CH=3 OP=3
cfg[4094] = { 1'b0, 8'hed, 8'h39}; // CH=1 OP=3
cfg[4095] = { 1'b0, 8'h79, 8'h53}; // CH=1 OP=2
cfg[4096] = { 1'b1, 8'h34, 8'hfb}; // CH=3 OP=1
cfg[4097] = { 1'b0, 8'hfc, 8'h63}; // CH=0 OP=3
cfg[4098] = { 1'b1, 8'hcd, 8'hcb}; // CH=4 OP=3
cfg[4099] = { 1'b0, 8'hb1, 8'hcc}; // CH=1 OP=0
cfg[4100] = { 1'b1, 8'hd9, 8'h55}; // CH=4 OP=2
cfg[4101] = { 1'b0, 8'hc9, 8'hf0}; // CH=1 OP=2
cfg[4102] = { 1'b0, 8'h6d, 8'hb6}; // CH=1 OP=3
cfg[4103] = { 1'b0, 8'hf6, 8'h45}; // CH=2 OP=1
cfg[4104] = { 1'b0, 8'he3, 8'h48}; // CH=3 OP=0
cfg[4105] = { 1'b0, 8'hd1, 8'h9b}; // CH=1 OP=0
cfg[4106] = { 1'b0, 8'h61, 8'hd}; // CH=1 OP=0
cfg[4107] = { 1'b0, 8'h5c, 8'h2}; // CH=0 OP=3
cfg[4108] = { 1'b1, 8'ha7, 8'hcf}; // CH=6 OP=1
cfg[4109] = { 1'b0, 8'hae, 8'h81}; // CH=2 OP=3
cfg[4110] = { 1'b1, 8'hd8, 8'h5a}; // CH=3 OP=2
cfg[4111] = { 1'b0, 8'h40, 8'h24}; // CH=0 OP=0
cfg[4112] = { 1'b0, 8'h49, 8'h91}; // CH=1 OP=2
cfg[4113] = { 1'b1, 8'h91, 8'h2a}; // CH=4 OP=0
cfg[4114] = { 1'b1, 8'h7d, 8'h83}; // CH=4 OP=3
cfg[4115] = { 1'b0, 8'h8a, 8'h27}; // CH=2 OP=2
cfg[4116] = { 1'b0, 8'hfa, 8'h88}; // CH=2 OP=2
cfg[4117] = { 1'b0, 8'h35, 8'he4}; // CH=1 OP=1
cfg[4118] = { 1'b0, 8'h3d, 8'h8b}; // CH=1 OP=3
cfg[4119] = { 1'b1, 8'h9b, 8'h39}; // CH=6 OP=2
cfg[4120] = { 1'b1, 8'he9, 8'h11}; // CH=4 OP=2
cfg[4121] = { 1'b1, 8'hed, 8'h51}; // CH=4 OP=3
cfg[4122] = { 1'b1, 8'h36, 8'h6a}; // CH=5 OP=1
cfg[4123] = { 1'b0, 8'hc8, 8'h94}; // CH=0 OP=2
cfg[4124] = { 1'b1, 8'hf4, 8'h17}; // CH=3 OP=1
cfg[4125] = { 1'b0, 8'hb6, 8'h6c}; // CH=2 OP=1
cfg[4126] = { 1'b0, 8'hb0, 8'ha3}; // CH=0 OP=0
cfg[4127] = { 1'b1, 8'he6, 8'h88}; // CH=5 OP=1
cfg[4128] = { 1'b1, 8'hfc, 8'h13}; // CH=3 OP=3
cfg[4129] = { 1'b1, 8'h5e, 8'hbe}; // CH=5 OP=3
cfg[4130] = { 1'b1, 8'hb0, 8'h2f}; // CH=3 OP=0
cfg[4131] = { 1'b0, 8'hcb, 8'hec}; // CH=3 OP=2
cfg[4132] = { 1'b0, 8'h93, 8'hae}; // CH=3 OP=0
cfg[4133] = { 1'b0, 8'h87, 8'hc6}; // CH=3 OP=1
cfg[4134] = { 1'b0, 8'ha3, 8'h32}; // CH=3 OP=0
cfg[4135] = { 1'b1, 8'h46, 8'hf8}; // CH=5 OP=1
cfg[4136] = { 1'b1, 8'hce, 8'h1b}; // CH=5 OP=3
cfg[4137] = { 1'b1, 8'he2, 8'h6a}; // CH=5 OP=0
cfg[4138] = { 1'b1, 8'h3b, 8'h66}; // CH=6 OP=2
cfg[4139] = { 1'b0, 8'he3, 8'h8d}; // CH=3 OP=0
cfg[4140] = { 1'b1, 8'h77, 8'h3d}; // CH=6 OP=1
cfg[4141] = { 1'b1, 8'h42, 8'h57}; // CH=5 OP=0
cfg[4142] = { 1'b1, 8'hd5, 8'h6}; // CH=4 OP=1
cfg[4143] = { 1'b1, 8'h5d, 8'hcc}; // CH=4 OP=3
cfg[4144] = { 1'b0, 8'h65, 8'hfe}; // CH=1 OP=1
cfg[4145] = { 1'b0, 8'hd8, 8'h46}; // CH=0 OP=2
cfg[4146] = { 1'b0, 8'h32, 8'h15}; // CH=2 OP=0
cfg[4147] = { 1'b0, 8'haf, 8'hf7}; // CH=3 OP=3
cfg[4148] = { 1'b1, 8'hea, 8'h26}; // CH=5 OP=2
cfg[4149] = { 1'b1, 8'hcd, 8'hb3}; // CH=4 OP=3
cfg[4150] = { 1'b0, 8'h45, 8'hf1}; // CH=1 OP=1
cfg[4151] = { 1'b1, 8'h87, 8'h48}; // CH=6 OP=1
cfg[4152] = { 1'b0, 8'h5d, 8'h4e}; // CH=1 OP=3
cfg[4153] = { 1'b0, 8'hba, 8'h1a}; // CH=2 OP=2
cfg[4154] = { 1'b0, 8'hba, 8'h18}; // CH=2 OP=2
cfg[4155] = { 1'b1, 8'h95, 8'hf}; // CH=4 OP=1
cfg[4156] = { 1'b1, 8'hc7, 8'h15}; // CH=6 OP=1
cfg[4157] = { 1'b1, 8'h76, 8'hc}; // CH=5 OP=1
cfg[4158] = { 1'b0, 8'h61, 8'h32}; // CH=1 OP=0
cfg[4159] = { 1'b1, 8'hb3, 8'he6}; // CH=6 OP=0
cfg[4160] = { 1'b1, 8'hfb, 8'h73}; // CH=6 OP=2
cfg[4161] = { 1'b1, 8'h58, 8'h6e}; // CH=3 OP=2
cfg[4162] = { 1'b1, 8'h4d, 8'h88}; // CH=4 OP=3
cfg[4163] = { 1'b1, 8'hb0, 8'hcc}; // CH=3 OP=0
cfg[4164] = { 1'b0, 8'hd1, 8'h9f}; // CH=1 OP=0
cfg[4165] = { 1'b0, 8'h6e, 8'h67}; // CH=2 OP=3
cfg[4166] = { 1'b0, 8'hef, 8'hdd}; // CH=3 OP=3
cfg[4167] = { 1'b1, 8'hbc, 8'h3e}; // CH=3 OP=3
cfg[4168] = { 1'b1, 8'h70, 8'h6d}; // CH=3 OP=0
cfg[4169] = { 1'b0, 8'h8e, 8'he0}; // CH=2 OP=3
cfg[4170] = { 1'b1, 8'hcd, 8'hdb}; // CH=4 OP=3
cfg[4171] = { 1'b1, 8'hc2, 8'h33}; // CH=5 OP=0
cfg[4172] = { 1'b0, 8'h95, 8'h45}; // CH=1 OP=1
cfg[4173] = { 1'b1, 8'h45, 8'h19}; // CH=4 OP=1
cfg[4174] = { 1'b0, 8'hc0, 8'hb9}; // CH=0 OP=0
cfg[4175] = { 1'b0, 8'hae, 8'h84}; // CH=2 OP=3
cfg[4176] = { 1'b1, 8'hcf, 8'h73}; // CH=6 OP=3
cfg[4177] = { 1'b0, 8'hd6, 8'h30}; // CH=2 OP=1
cfg[4178] = { 1'b1, 8'hb4, 8'ha0}; // CH=3 OP=1
cfg[4179] = { 1'b1, 8'hb2, 8'h2e}; // CH=5 OP=0
cfg[4180] = { 1'b1, 8'h98, 8'hfc}; // CH=3 OP=2
cfg[4181] = { 1'b0, 8'hde, 8'h11}; // CH=2 OP=3
cfg[4182] = { 1'b0, 8'hef, 8'ha6}; // CH=3 OP=3
cfg[4183] = { 1'b1, 8'hcd, 8'heb}; // CH=4 OP=3
cfg[4184] = { 1'b0, 8'h8d, 8'h1}; // CH=1 OP=3
cfg[4185] = { 1'b0, 8'h3c, 8'h86}; // CH=0 OP=3
cfg[4186] = { 1'b0, 8'hfa, 8'hf9}; // CH=2 OP=2
cfg[4187] = { 1'b1, 8'ha3, 8'he2}; // CH=6 OP=0
cfg[4188] = { 1'b1, 8'hf8, 8'h96}; // CH=3 OP=2
cfg[4189] = { 1'b0, 8'hf4, 8'h91}; // CH=0 OP=1
cfg[4190] = { 1'b0, 8'hb2, 8'h2a}; // CH=2 OP=0
cfg[4191] = { 1'b1, 8'h80, 8'h8}; // CH=3 OP=0
cfg[4192] = { 1'b0, 8'h68, 8'hf7}; // CH=0 OP=2
cfg[4193] = { 1'b1, 8'h52, 8'hc5}; // CH=5 OP=0
cfg[4194] = { 1'b1, 8'h8e, 8'h91}; // CH=5 OP=3
cfg[4195] = { 1'b1, 8'h9a, 8'h8a}; // CH=5 OP=2
cfg[4196] = { 1'b1, 8'h7c, 8'hb4}; // CH=3 OP=3
cfg[4197] = { 1'b0, 8'h50, 8'h7d}; // CH=0 OP=0
cfg[4198] = { 1'b1, 8'he2, 8'h5b}; // CH=5 OP=0
cfg[4199] = { 1'b1, 8'h38, 8'hc1}; // CH=3 OP=2
cfg[4200] = { 1'b0, 8'h56, 8'h9c}; // CH=2 OP=1
cfg[4201] = { 1'b1, 8'h60, 8'h4}; // CH=3 OP=0
cfg[4202] = { 1'b0, 8'h6b, 8'hd}; // CH=3 OP=2
cfg[4203] = { 1'b1, 8'hfc, 8'hd6}; // CH=3 OP=3
cfg[4204] = { 1'b1, 8'h86, 8'h5d}; // CH=5 OP=1
cfg[4205] = { 1'b1, 8'h3a, 8'hde}; // CH=5 OP=2
cfg[4206] = { 1'b1, 8'hb8, 8'h2}; // CH=3 OP=2
cfg[4207] = { 1'b0, 8'h35, 8'h52}; // CH=1 OP=1
cfg[4208] = { 1'b0, 8'hf6, 8'h97}; // CH=2 OP=1
cfg[4209] = { 1'b0, 8'h54, 8'hb3}; // CH=0 OP=1
cfg[4210] = { 1'b1, 8'h60, 8'h85}; // CH=3 OP=0
cfg[4211] = { 1'b0, 8'h30, 8'he5}; // CH=0 OP=0
cfg[4212] = { 1'b1, 8'h53, 8'h50}; // CH=6 OP=0
cfg[4213] = { 1'b1, 8'h94, 8'h4c}; // CH=3 OP=1
cfg[4214] = { 1'b0, 8'h72, 8'h50}; // CH=2 OP=0
cfg[4215] = { 1'b1, 8'h74, 8'h18}; // CH=3 OP=1
cfg[4216] = { 1'b1, 8'hc6, 8'hf2}; // CH=5 OP=1
cfg[4217] = { 1'b0, 8'hfb, 8'h27}; // CH=3 OP=2
cfg[4218] = { 1'b1, 8'h3b, 8'h1d}; // CH=6 OP=2
cfg[4219] = { 1'b0, 8'h90, 8'h4b}; // CH=0 OP=0
cfg[4220] = { 1'b0, 8'hf0, 8'hd0}; // CH=0 OP=0
cfg[4221] = { 1'b0, 8'h41, 8'hb5}; // CH=1 OP=0
cfg[4222] = { 1'b1, 8'h78, 8'h74}; // CH=3 OP=2
cfg[4223] = { 1'b1, 8'hc9, 8'h79}; // CH=4 OP=2
cfg[4224] = { 1'b0, 8'he1, 8'h31}; // CH=1 OP=0
cfg[4225] = { 1'b0, 8'hd3, 8'hf6}; // CH=3 OP=0
cfg[4226] = { 1'b0, 8'hfa, 8'he8}; // CH=2 OP=2
cfg[4227] = { 1'b1, 8'hef, 8'h72}; // CH=6 OP=3
cfg[4228] = { 1'b0, 8'h7f, 8'h63}; // CH=3 OP=3
cfg[4229] = { 1'b0, 8'h6f, 8'h33}; // CH=3 OP=3
cfg[4230] = { 1'b0, 8'h8f, 8'he9}; // CH=3 OP=3
cfg[4231] = { 1'b1, 8'hd3, 8'hee}; // CH=6 OP=0
cfg[4232] = { 1'b0, 8'hdf, 8'h7c}; // CH=3 OP=3
cfg[4233] = { 1'b0, 8'h5d, 8'h46}; // CH=1 OP=3
cfg[4234] = { 1'b1, 8'h4f, 8'h27}; // CH=6 OP=3
cfg[4235] = { 1'b1, 8'h73, 8'hfb}; // CH=6 OP=0
cfg[4236] = { 1'b1, 8'he5, 8'hbb}; // CH=4 OP=1
cfg[4237] = { 1'b1, 8'h94, 8'haa}; // CH=3 OP=1
cfg[4238] = { 1'b0, 8'hce, 8'h29}; // CH=2 OP=3
cfg[4239] = { 1'b1, 8'he9, 8'h98}; // CH=4 OP=2
cfg[4240] = { 1'b0, 8'h44, 8'h28}; // CH=0 OP=1
cfg[4241] = { 1'b1, 8'hbb, 8'h2b}; // CH=6 OP=2
cfg[4242] = { 1'b0, 8'hee, 8'hf7}; // CH=2 OP=3
cfg[4243] = { 1'b1, 8'ha4, 8'hb4}; // CH=3 OP=1
cfg[4244] = { 1'b1, 8'hac, 8'h10}; // CH=3 OP=3
cfg[4245] = { 1'b0, 8'h68, 8'h6}; // CH=0 OP=2
cfg[4246] = { 1'b0, 8'h83, 8'h13}; // CH=3 OP=0
cfg[4247] = { 1'b0, 8'hd4, 8'hfa}; // CH=0 OP=1
cfg[4248] = { 1'b1, 8'hfc, 8'hb3}; // CH=3 OP=3
cfg[4249] = { 1'b0, 8'h40, 8'h2e}; // CH=0 OP=0
cfg[4250] = { 1'b1, 8'h37, 8'hd0}; // CH=6 OP=1
cfg[4251] = { 1'b0, 8'h8c, 8'hbe}; // CH=0 OP=3
cfg[4252] = { 1'b0, 8'h31, 8'hd3}; // CH=1 OP=0
cfg[4253] = { 1'b1, 8'hdd, 8'he4}; // CH=4 OP=3
cfg[4254] = { 1'b1, 8'h45, 8'hea}; // CH=4 OP=1
cfg[4255] = { 1'b1, 8'h58, 8'hfd}; // CH=3 OP=2
cfg[4256] = { 1'b1, 8'h94, 8'h80}; // CH=3 OP=1
cfg[4257] = { 1'b0, 8'h68, 8'ha6}; // CH=0 OP=2
cfg[4258] = { 1'b1, 8'h65, 8'h59}; // CH=4 OP=1
cfg[4259] = { 1'b1, 8'h8d, 8'h87}; // CH=4 OP=3
cfg[4260] = { 1'b1, 8'h5d, 8'h70}; // CH=4 OP=3
cfg[4261] = { 1'b1, 8'h7b, 8'h78}; // CH=6 OP=2
cfg[4262] = { 1'b0, 8'hac, 8'hee}; // CH=0 OP=3
cfg[4263] = { 1'b1, 8'h8a, 8'hd2}; // CH=5 OP=2
cfg[4264] = { 1'b1, 8'hcf, 8'hbc}; // CH=6 OP=3
cfg[4265] = { 1'b0, 8'h94, 8'hb9}; // CH=0 OP=1
cfg[4266] = { 1'b1, 8'he0, 8'hbb}; // CH=3 OP=0
cfg[4267] = { 1'b0, 8'h39, 8'h4f}; // CH=1 OP=2
cfg[4268] = { 1'b1, 8'hc1, 8'hc7}; // CH=4 OP=0
cfg[4269] = { 1'b0, 8'h31, 8'h7e}; // CH=1 OP=0
cfg[4270] = { 1'b1, 8'haa, 8'h6d}; // CH=5 OP=2
cfg[4271] = { 1'b0, 8'hde, 8'he9}; // CH=2 OP=3
cfg[4272] = { 1'b0, 8'h4f, 8'h95}; // CH=3 OP=3
cfg[4273] = { 1'b1, 8'hef, 8'heb}; // CH=6 OP=3
cfg[4274] = { 1'b1, 8'ha1, 8'hc5}; // CH=4 OP=0
cfg[4275] = { 1'b0, 8'ha1, 8'hd2}; // CH=1 OP=0
cfg[4276] = { 1'b0, 8'hf1, 8'hf6}; // CH=1 OP=0
cfg[4277] = { 1'b0, 8'hb8, 8'h7f}; // CH=0 OP=2
cfg[4278] = { 1'b1, 8'h36, 8'h95}; // CH=5 OP=1
cfg[4279] = { 1'b0, 8'ha4, 8'h8}; // CH=0 OP=1
cfg[4280] = { 1'b0, 8'h8d, 8'h96}; // CH=1 OP=3
cfg[4281] = { 1'b1, 8'ha1, 8'h12}; // CH=4 OP=0
cfg[4282] = { 1'b1, 8'h8c, 8'h42}; // CH=3 OP=3
cfg[4283] = { 1'b1, 8'h99, 8'h31}; // CH=4 OP=2
cfg[4284] = { 1'b0, 8'h3b, 8'h47}; // CH=3 OP=2
cfg[4285] = { 1'b0, 8'hdc, 8'h19}; // CH=0 OP=3
cfg[4286] = { 1'b1, 8'hcd, 8'hf}; // CH=4 OP=3
cfg[4287] = { 1'b1, 8'h85, 8'h8e}; // CH=4 OP=1
cfg[4288] = { 1'b0, 8'hbc, 8'h23}; // CH=0 OP=3
cfg[4289] = { 1'b0, 8'h60, 8'h2b}; // CH=0 OP=0
cfg[4290] = { 1'b1, 8'hed, 8'hc1}; // CH=4 OP=3
cfg[4291] = { 1'b0, 8'hf3, 8'hd4}; // CH=3 OP=0
cfg[4292] = { 1'b1, 8'h7f, 8'h51}; // CH=6 OP=3
cfg[4293] = { 1'b0, 8'hd4, 8'h82}; // CH=0 OP=1
cfg[4294] = { 1'b0, 8'he3, 8'h53}; // CH=3 OP=0
cfg[4295] = { 1'b0, 8'hf3, 8'h14}; // CH=3 OP=0
cfg[4296] = { 1'b1, 8'h81, 8'h3b}; // CH=4 OP=0
cfg[4297] = { 1'b1, 8'ha5, 8'h3b}; // CH=4 OP=1
cfg[4298] = { 1'b1, 8'hd0, 8'h45}; // CH=3 OP=0
cfg[4299] = { 1'b1, 8'h92, 8'h4}; // CH=5 OP=0
cfg[4300] = { 1'b0, 8'h66, 8'h56}; // CH=2 OP=1
cfg[4301] = { 1'b1, 8'h9b, 8'h49}; // CH=6 OP=2
cfg[4302] = { 1'b1, 8'h3e, 8'hc8}; // CH=5 OP=3
cfg[4303] = { 1'b1, 8'h39, 8'he1}; // CH=4 OP=2
cfg[4304] = { 1'b0, 8'h64, 8'h17}; // CH=0 OP=1
cfg[4305] = { 1'b1, 8'h62, 8'h10}; // CH=5 OP=0
cfg[4306] = { 1'b0, 8'he5, 8'h91}; // CH=1 OP=1
cfg[4307] = { 1'b1, 8'he7, 8'h36}; // CH=6 OP=1
cfg[4308] = { 1'b1, 8'heb, 8'hc3}; // CH=6 OP=2
cfg[4309] = { 1'b1, 8'h42, 8'h4f}; // CH=5 OP=0
cfg[4310] = { 1'b1, 8'h8b, 8'hea}; // CH=6 OP=2
cfg[4311] = { 1'b0, 8'h54, 8'hd7}; // CH=0 OP=1
cfg[4312] = { 1'b0, 8'h35, 8'h47}; // CH=1 OP=1
cfg[4313] = { 1'b1, 8'h69, 8'h80}; // CH=4 OP=2
cfg[4314] = { 1'b0, 8'hce, 8'h9d}; // CH=2 OP=3
cfg[4315] = { 1'b0, 8'h30, 8'had}; // CH=0 OP=0
cfg[4316] = { 1'b0, 8'h36, 8'h3f}; // CH=2 OP=1
cfg[4317] = { 1'b1, 8'h7c, 8'h39}; // CH=3 OP=3
cfg[4318] = { 1'b0, 8'h4b, 8'h8}; // CH=3 OP=2
cfg[4319] = { 1'b0, 8'h35, 8'h14}; // CH=1 OP=1
cfg[4320] = { 1'b0, 8'h87, 8'haf}; // CH=3 OP=1
cfg[4321] = { 1'b0, 8'h72, 8'h5f}; // CH=2 OP=0
cfg[4322] = { 1'b0, 8'h75, 8'hc8}; // CH=1 OP=1
cfg[4323] = { 1'b0, 8'ha3, 8'h96}; // CH=3 OP=0
cfg[4324] = { 1'b1, 8'h37, 8'hc6}; // CH=6 OP=1
cfg[4325] = { 1'b0, 8'h6d, 8'hdb}; // CH=1 OP=3
cfg[4326] = { 1'b0, 8'h8a, 8'h14}; // CH=2 OP=2
cfg[4327] = { 1'b0, 8'h93, 8'h10}; // CH=3 OP=0
cfg[4328] = { 1'b0, 8'hdd, 8'h5b}; // CH=1 OP=3
cfg[4329] = { 1'b0, 8'hb3, 8'h91}; // CH=3 OP=0
cfg[4330] = { 1'b1, 8'hdd, 8'h9e}; // CH=4 OP=3
cfg[4331] = { 1'b1, 8'h3c, 8'hf2}; // CH=3 OP=3
cfg[4332] = { 1'b1, 8'h98, 8'hc6}; // CH=3 OP=2
cfg[4333] = { 1'b0, 8'h3b, 8'h9b}; // CH=3 OP=2
cfg[4334] = { 1'b0, 8'h73, 8'h62}; // CH=3 OP=0
cfg[4335] = { 1'b0, 8'he0, 8'h3d}; // CH=0 OP=0
cfg[4336] = { 1'b0, 8'h6b, 8'h52}; // CH=3 OP=2
cfg[4337] = { 1'b1, 8'hfe, 8'h62}; // CH=5 OP=3
cfg[4338] = { 1'b1, 8'hdb, 8'hbe}; // CH=6 OP=2
cfg[4339] = { 1'b1, 8'h8f, 8'h4f}; // CH=6 OP=3
cfg[4340] = { 1'b1, 8'h6c, 8'hed}; // CH=3 OP=3
cfg[4341] = { 1'b0, 8'ha9, 8'hdf}; // CH=1 OP=2
cfg[4342] = { 1'b1, 8'hae, 8'ha5}; // CH=5 OP=3
cfg[4343] = { 1'b0, 8'h49, 8'hde}; // CH=1 OP=2
cfg[4344] = { 1'b1, 8'hab, 8'h36}; // CH=6 OP=2
cfg[4345] = { 1'b0, 8'he9, 8'hec}; // CH=1 OP=2
cfg[4346] = { 1'b1, 8'h3b, 8'h77}; // CH=6 OP=2
cfg[4347] = { 1'b0, 8'h9d, 8'h52}; // CH=1 OP=3
cfg[4348] = { 1'b0, 8'h5b, 8'h93}; // CH=3 OP=2
cfg[4349] = { 1'b1, 8'haa, 8'h4e}; // CH=5 OP=2
cfg[4350] = { 1'b0, 8'h97, 8'h33}; // CH=3 OP=1
cfg[4351] = { 1'b1, 8'h76, 8'hc9}; // CH=5 OP=1
cfg[4352] = { 1'b0, 8'h78, 8'h83}; // CH=0 OP=2
cfg[4353] = { 1'b1, 8'hc1, 8'hfa}; // CH=4 OP=0
cfg[4354] = { 1'b0, 8'h6d, 8'h30}; // CH=1 OP=3
cfg[4355] = { 1'b1, 8'h56, 8'h1c}; // CH=5 OP=1
cfg[4356] = { 1'b0, 8'h91, 8'h93}; // CH=1 OP=0
cfg[4357] = { 1'b0, 8'hda, 8'he5}; // CH=2 OP=2
cfg[4358] = { 1'b0, 8'hff, 8'h8a}; // CH=3 OP=3
cfg[4359] = { 1'b1, 8'hb4, 8'h34}; // CH=3 OP=1
cfg[4360] = { 1'b0, 8'hd5, 8'hcc}; // CH=1 OP=1
cfg[4361] = { 1'b0, 8'h9f, 8'h42}; // CH=3 OP=3
cfg[4362] = { 1'b1, 8'h58, 8'h5e}; // CH=3 OP=2
cfg[4363] = { 1'b0, 8'h88, 8'h7e}; // CH=0 OP=2
cfg[4364] = { 1'b1, 8'ha5, 8'he1}; // CH=4 OP=1
cfg[4365] = { 1'b1, 8'h38, 8'h25}; // CH=3 OP=2
cfg[4366] = { 1'b0, 8'h5b, 8'hb5}; // CH=3 OP=2
cfg[4367] = { 1'b1, 8'he5, 8'h96}; // CH=4 OP=1
cfg[4368] = { 1'b1, 8'h43, 8'h5d}; // CH=6 OP=0
cfg[4369] = { 1'b0, 8'hb7, 8'he5}; // CH=3 OP=1
cfg[4370] = { 1'b1, 8'hce, 8'h86}; // CH=5 OP=3
cfg[4371] = { 1'b1, 8'ha6, 8'hdf}; // CH=5 OP=1
cfg[4372] = { 1'b1, 8'hec, 8'h67}; // CH=3 OP=3
cfg[4373] = { 1'b1, 8'h87, 8'hc}; // CH=6 OP=1
cfg[4374] = { 1'b0, 8'hb4, 8'h45}; // CH=0 OP=1
cfg[4375] = { 1'b0, 8'h49, 8'h63}; // CH=1 OP=2
cfg[4376] = { 1'b1, 8'hd8, 8'hf4}; // CH=3 OP=2
cfg[4377] = { 1'b1, 8'haf, 8'hd}; // CH=6 OP=3
cfg[4378] = { 1'b1, 8'hcb, 8'h33}; // CH=6 OP=2
cfg[4379] = { 1'b1, 8'ha1, 8'hea}; // CH=4 OP=0
cfg[4380] = { 1'b0, 8'h80, 8'had}; // CH=0 OP=0
cfg[4381] = { 1'b1, 8'he8, 8'haa}; // CH=3 OP=2
cfg[4382] = { 1'b1, 8'hf4, 8'h89}; // CH=3 OP=1
cfg[4383] = { 1'b0, 8'h39, 8'h8e}; // CH=1 OP=2
cfg[4384] = { 1'b0, 8'h9c, 8'h48}; // CH=0 OP=3
cfg[4385] = { 1'b1, 8'h96, 8'h91}; // CH=5 OP=1
cfg[4386] = { 1'b1, 8'hed, 8'h6a}; // CH=4 OP=3
cfg[4387] = { 1'b1, 8'h9c, 8'h85}; // CH=3 OP=3
cfg[4388] = { 1'b0, 8'h67, 8'hb9}; // CH=3 OP=1
cfg[4389] = { 1'b1, 8'h95, 8'ha3}; // CH=4 OP=1
cfg[4390] = { 1'b0, 8'h42, 8'h5c}; // CH=2 OP=0
cfg[4391] = { 1'b1, 8'hec, 8'hbb}; // CH=3 OP=3
cfg[4392] = { 1'b1, 8'h76, 8'h6}; // CH=5 OP=1
cfg[4393] = { 1'b1, 8'hdd, 8'hd8}; // CH=4 OP=3
cfg[4394] = { 1'b1, 8'h79, 8'h4c}; // CH=4 OP=2
cfg[4395] = { 1'b0, 8'h7e, 8'hdd}; // CH=2 OP=3
cfg[4396] = { 1'b1, 8'hcd, 8'hfc}; // CH=4 OP=3
cfg[4397] = { 1'b0, 8'h86, 8'h9f}; // CH=2 OP=1
cfg[4398] = { 1'b1, 8'h94, 8'h44}; // CH=3 OP=1
cfg[4399] = { 1'b0, 8'hd6, 8'h85}; // CH=2 OP=1
cfg[4400] = { 1'b1, 8'hc3, 8'h40}; // CH=6 OP=0
cfg[4401] = { 1'b0, 8'h39, 8'h46}; // CH=1 OP=2
cfg[4402] = { 1'b0, 8'h3d, 8'h1f}; // CH=1 OP=3
cfg[4403] = { 1'b1, 8'h89, 8'h7e}; // CH=4 OP=2
cfg[4404] = { 1'b0, 8'h66, 8'h72}; // CH=2 OP=1
cfg[4405] = { 1'b0, 8'hae, 8'hf0}; // CH=2 OP=3
cfg[4406] = { 1'b0, 8'h7b, 8'h5}; // CH=3 OP=2
cfg[4407] = { 1'b1, 8'h9e, 8'ha4}; // CH=5 OP=3
cfg[4408] = { 1'b0, 8'h33, 8'h2a}; // CH=3 OP=0
cfg[4409] = { 1'b1, 8'hc4, 8'hb0}; // CH=3 OP=1
cfg[4410] = { 1'b0, 8'hc5, 8'hcc}; // CH=1 OP=1
cfg[4411] = { 1'b1, 8'h69, 8'h5}; // CH=4 OP=2
cfg[4412] = { 1'b0, 8'hea, 8'h42}; // CH=2 OP=2
cfg[4413] = { 1'b0, 8'he4, 8'hcb}; // CH=0 OP=1
cfg[4414] = { 1'b0, 8'hee, 8'h32}; // CH=2 OP=3
cfg[4415] = { 1'b1, 8'hf5, 8'he0}; // CH=4 OP=1
cfg[4416] = { 1'b0, 8'h94, 8'h5b}; // CH=0 OP=1
cfg[4417] = { 1'b1, 8'h32, 8'h5c}; // CH=5 OP=0
cfg[4418] = { 1'b1, 8'h65, 8'h86}; // CH=4 OP=1
cfg[4419] = { 1'b0, 8'h6f, 8'h36}; // CH=3 OP=3
cfg[4420] = { 1'b1, 8'h3b, 8'h27}; // CH=6 OP=2
cfg[4421] = { 1'b0, 8'h41, 8'h5e}; // CH=1 OP=0
cfg[4422] = { 1'b1, 8'h83, 8'hb4}; // CH=6 OP=0
cfg[4423] = { 1'b1, 8'h4f, 8'h88}; // CH=6 OP=3
cfg[4424] = { 1'b1, 8'h81, 8'hce}; // CH=4 OP=0
cfg[4425] = { 1'b0, 8'h61, 8'h5}; // CH=1 OP=0
cfg[4426] = { 1'b1, 8'hbc, 8'h42}; // CH=3 OP=3
cfg[4427] = { 1'b1, 8'ha7, 8'h23}; // CH=6 OP=1
cfg[4428] = { 1'b0, 8'hd5, 8'h9e}; // CH=1 OP=1
cfg[4429] = { 1'b0, 8'hfc, 8'h2a}; // CH=0 OP=3
cfg[4430] = { 1'b1, 8'h5a, 8'hf0}; // CH=5 OP=2
cfg[4431] = { 1'b0, 8'h7c, 8'h1f}; // CH=0 OP=3
cfg[4432] = { 1'b0, 8'hcb, 8'h96}; // CH=3 OP=2
cfg[4433] = { 1'b1, 8'h4c, 8'h64}; // CH=3 OP=3
cfg[4434] = { 1'b1, 8'had, 8'h6a}; // CH=4 OP=3
cfg[4435] = { 1'b0, 8'h69, 8'hac}; // CH=1 OP=2
cfg[4436] = { 1'b1, 8'h81, 8'hcf}; // CH=4 OP=0
cfg[4437] = { 1'b1, 8'he4, 8'hbb}; // CH=3 OP=1
cfg[4438] = { 1'b0, 8'hf0, 8'ha8}; // CH=0 OP=0
cfg[4439] = { 1'b1, 8'h4a, 8'hfe}; // CH=5 OP=2
cfg[4440] = { 1'b0, 8'h58, 8'h1d}; // CH=0 OP=2
cfg[4441] = { 1'b0, 8'hee, 8'h55}; // CH=2 OP=3
cfg[4442] = { 1'b1, 8'h53, 8'h8b}; // CH=6 OP=0
cfg[4443] = { 1'b1, 8'hbd, 8'hac}; // CH=4 OP=3
cfg[4444] = { 1'b0, 8'h69, 8'haf}; // CH=1 OP=2
cfg[4445] = { 1'b1, 8'h38, 8'h26}; // CH=3 OP=2
cfg[4446] = { 1'b0, 8'hf3, 8'h45}; // CH=3 OP=0
cfg[4447] = { 1'b1, 8'hd8, 8'h71}; // CH=3 OP=2
cfg[4448] = { 1'b0, 8'he6, 8'h19}; // CH=2 OP=1
cfg[4449] = { 1'b0, 8'he5, 8'h79}; // CH=1 OP=1
cfg[4450] = { 1'b1, 8'ha5, 8'hd1}; // CH=4 OP=1
cfg[4451] = { 1'b0, 8'h44, 8'h18}; // CH=0 OP=1
cfg[4452] = { 1'b1, 8'h8f, 8'h6b}; // CH=6 OP=3
cfg[4453] = { 1'b0, 8'h3e, 8'hc7}; // CH=2 OP=3
cfg[4454] = { 1'b1, 8'h65, 8'hc8}; // CH=4 OP=1
cfg[4455] = { 1'b1, 8'haa, 8'h4a}; // CH=5 OP=2
cfg[4456] = { 1'b0, 8'h94, 8'heb}; // CH=0 OP=1
cfg[4457] = { 1'b1, 8'h7b, 8'h35}; // CH=6 OP=2
cfg[4458] = { 1'b0, 8'h60, 8'hae}; // CH=0 OP=0
cfg[4459] = { 1'b1, 8'h62, 8'h7f}; // CH=5 OP=0
cfg[4460] = { 1'b0, 8'hba, 8'h24}; // CH=2 OP=2
cfg[4461] = { 1'b0, 8'h9d, 8'h68}; // CH=1 OP=3
cfg[4462] = { 1'b1, 8'had, 8'h97}; // CH=4 OP=3
cfg[4463] = { 1'b0, 8'h3e, 8'h6b}; // CH=2 OP=3
cfg[4464] = { 1'b0, 8'h70, 8'hd0}; // CH=0 OP=0
cfg[4465] = { 1'b1, 8'h5c, 8'hc4}; // CH=3 OP=3
cfg[4466] = { 1'b1, 8'hdd, 8'h58}; // CH=4 OP=3
cfg[4467] = { 1'b0, 8'he5, 8'hd3}; // CH=1 OP=1
cfg[4468] = { 1'b1, 8'hbe, 8'h33}; // CH=5 OP=3
cfg[4469] = { 1'b0, 8'hc1, 8'h96}; // CH=1 OP=0
cfg[4470] = { 1'b1, 8'hdb, 8'h50}; // CH=6 OP=2
cfg[4471] = { 1'b1, 8'h61, 8'hee}; // CH=4 OP=0
cfg[4472] = { 1'b1, 8'h7d, 8'h1b}; // CH=4 OP=3
cfg[4473] = { 1'b0, 8'ha4, 8'h4d}; // CH=0 OP=1
cfg[4474] = { 1'b1, 8'hd2, 8'h54}; // CH=5 OP=0
cfg[4475] = { 1'b0, 8'h69, 8'h70}; // CH=1 OP=2
cfg[4476] = { 1'b1, 8'h35, 8'h4e}; // CH=4 OP=1
cfg[4477] = { 1'b0, 8'hb0, 8'h33}; // CH=0 OP=0
cfg[4478] = { 1'b0, 8'hab, 8'hf2}; // CH=3 OP=2
cfg[4479] = { 1'b0, 8'hca, 8'hb3}; // CH=2 OP=2
cfg[4480] = { 1'b0, 8'h51, 8'h8e}; // CH=1 OP=0
cfg[4481] = { 1'b0, 8'h70, 8'hef}; // CH=0 OP=0
cfg[4482] = { 1'b1, 8'hee, 8'hfe}; // CH=5 OP=3
cfg[4483] = { 1'b0, 8'h92, 8'h4b}; // CH=2 OP=0
cfg[4484] = { 1'b1, 8'ha6, 8'h9f}; // CH=5 OP=1
cfg[4485] = { 1'b1, 8'h80, 8'hb8}; // CH=3 OP=0
cfg[4486] = { 1'b1, 8'hb5, 8'h65}; // CH=4 OP=1
cfg[4487] = { 1'b1, 8'h66, 8'h98}; // CH=5 OP=1
cfg[4488] = { 1'b1, 8'hf3, 8'h8a}; // CH=6 OP=0
cfg[4489] = { 1'b1, 8'h52, 8'hdb}; // CH=5 OP=0
cfg[4490] = { 1'b0, 8'h9e, 8'h2c}; // CH=2 OP=3
cfg[4491] = { 1'b1, 8'hb9, 8'h9d}; // CH=4 OP=2
cfg[4492] = { 1'b1, 8'h39, 8'hf4}; // CH=4 OP=2
cfg[4493] = { 1'b0, 8'h50, 8'hc3}; // CH=0 OP=0
cfg[4494] = { 1'b0, 8'hd0, 8'hda}; // CH=0 OP=0
cfg[4495] = { 1'b1, 8'h85, 8'h3f}; // CH=4 OP=1
cfg[4496] = { 1'b0, 8'heb, 8'hd8}; // CH=3 OP=2
cfg[4497] = { 1'b0, 8'hfc, 8'h62}; // CH=0 OP=3
cfg[4498] = { 1'b1, 8'hd7, 8'ha0}; // CH=6 OP=1
cfg[4499] = { 1'b1, 8'hbc, 8'h6c}; // CH=3 OP=3
cfg[4500] = { 1'b1, 8'hc2, 8'ha1}; // CH=5 OP=0
cfg[4501] = { 1'b1, 8'hb6, 8'h2c}; // CH=5 OP=1
cfg[4502] = { 1'b1, 8'hef, 8'h49}; // CH=6 OP=3
cfg[4503] = { 1'b1, 8'h3f, 8'hc}; // CH=6 OP=3
cfg[4504] = { 1'b1, 8'h6a, 8'he7}; // CH=5 OP=2
cfg[4505] = { 1'b0, 8'h5d, 8'h94}; // CH=1 OP=3
cfg[4506] = { 1'b0, 8'h35, 8'h80}; // CH=1 OP=1
cfg[4507] = { 1'b1, 8'h54, 8'h7c}; // CH=3 OP=1
cfg[4508] = { 1'b0, 8'h58, 8'h6d}; // CH=0 OP=2
cfg[4509] = { 1'b0, 8'hf9, 8'h94}; // CH=1 OP=2
cfg[4510] = { 1'b0, 8'h52, 8'h75}; // CH=2 OP=0
cfg[4511] = { 1'b1, 8'h41, 8'h6e}; // CH=4 OP=0
cfg[4512] = { 1'b0, 8'h80, 8'h7a}; // CH=0 OP=0
cfg[4513] = { 1'b0, 8'h8f, 8'h61}; // CH=3 OP=3
cfg[4514] = { 1'b0, 8'h91, 8'h88}; // CH=1 OP=0
cfg[4515] = { 1'b0, 8'hc6, 8'ha3}; // CH=2 OP=1
cfg[4516] = { 1'b1, 8'hc7, 8'h20}; // CH=6 OP=1
cfg[4517] = { 1'b0, 8'he5, 8'h74}; // CH=1 OP=1
cfg[4518] = { 1'b1, 8'hbf, 8'hcc}; // CH=6 OP=3
cfg[4519] = { 1'b0, 8'h5b, 8'hc5}; // CH=3 OP=2
cfg[4520] = { 1'b1, 8'had, 8'hea}; // CH=4 OP=3
cfg[4521] = { 1'b0, 8'hee, 8'h58}; // CH=2 OP=3
cfg[4522] = { 1'b1, 8'h6e, 8'hd2}; // CH=5 OP=3
cfg[4523] = { 1'b1, 8'hfd, 8'h34}; // CH=4 OP=3
cfg[4524] = { 1'b1, 8'h42, 8'hbc}; // CH=5 OP=0
cfg[4525] = { 1'b0, 8'he4, 8'hf5}; // CH=0 OP=1
cfg[4526] = { 1'b0, 8'h58, 8'h12}; // CH=0 OP=2
cfg[4527] = { 1'b1, 8'h60, 8'h68}; // CH=3 OP=0
cfg[4528] = { 1'b0, 8'hbb, 8'he9}; // CH=3 OP=2
cfg[4529] = { 1'b1, 8'h68, 8'hd3}; // CH=3 OP=2
cfg[4530] = { 1'b0, 8'h56, 8'h2b}; // CH=2 OP=1
cfg[4531] = { 1'b1, 8'hc4, 8'hfd}; // CH=3 OP=1
cfg[4532] = { 1'b0, 8'hc1, 8'h31}; // CH=1 OP=0
cfg[4533] = { 1'b1, 8'he2, 8'hed}; // CH=5 OP=0
cfg[4534] = { 1'b0, 8'ha6, 8'h30}; // CH=2 OP=1
cfg[4535] = { 1'b0, 8'h8a, 8'h5a}; // CH=2 OP=2
cfg[4536] = { 1'b0, 8'he2, 8'h6c}; // CH=2 OP=0
cfg[4537] = { 1'b0, 8'hf4, 8'hd4}; // CH=0 OP=1
cfg[4538] = { 1'b0, 8'hb0, 8'hef}; // CH=0 OP=0
cfg[4539] = { 1'b0, 8'h44, 8'hc2}; // CH=0 OP=1
cfg[4540] = { 1'b1, 8'h4f, 8'h6f}; // CH=6 OP=3
cfg[4541] = { 1'b0, 8'hc3, 8'h33}; // CH=3 OP=0
cfg[4542] = { 1'b0, 8'hd4, 8'hf5}; // CH=0 OP=1
cfg[4543] = { 1'b1, 8'h39, 8'hd7}; // CH=4 OP=2
cfg[4544] = { 1'b1, 8'h93, 8'h4b}; // CH=6 OP=0
cfg[4545] = { 1'b1, 8'he9, 8'h3d}; // CH=4 OP=2
cfg[4546] = { 1'b1, 8'hef, 8'hd4}; // CH=6 OP=3
cfg[4547] = { 1'b0, 8'hde, 8'hfb}; // CH=2 OP=3
cfg[4548] = { 1'b0, 8'ha0, 8'hd3}; // CH=0 OP=0
cfg[4549] = { 1'b0, 8'h8d, 8'h17}; // CH=1 OP=3
cfg[4550] = { 1'b1, 8'h77, 8'h66}; // CH=6 OP=1
cfg[4551] = { 1'b1, 8'h93, 8'h29}; // CH=6 OP=0
cfg[4552] = { 1'b0, 8'h9d, 8'hfd}; // CH=1 OP=3
cfg[4553] = { 1'b1, 8'hd6, 8'h12}; // CH=5 OP=1
cfg[4554] = { 1'b0, 8'h6a, 8'h5d}; // CH=2 OP=2
cfg[4555] = { 1'b1, 8'h6a, 8'h9b}; // CH=5 OP=2
cfg[4556] = { 1'b0, 8'h3e, 8'h6c}; // CH=2 OP=3
cfg[4557] = { 1'b1, 8'h39, 8'h32}; // CH=4 OP=2
cfg[4558] = { 1'b1, 8'hd7, 8'ha8}; // CH=6 OP=1
cfg[4559] = { 1'b1, 8'h64, 8'h23}; // CH=3 OP=1
cfg[4560] = { 1'b0, 8'hdb, 8'h89}; // CH=3 OP=2
cfg[4561] = { 1'b1, 8'h6f, 8'hb2}; // CH=6 OP=3
cfg[4562] = { 1'b1, 8'h88, 8'hb0}; // CH=3 OP=2
cfg[4563] = { 1'b0, 8'h4c, 8'he2}; // CH=0 OP=3
cfg[4564] = { 1'b1, 8'hb6, 8'hbb}; // CH=5 OP=1
cfg[4565] = { 1'b1, 8'hf5, 8'h27}; // CH=4 OP=1
cfg[4566] = { 1'b0, 8'h7d, 8'h5a}; // CH=1 OP=3
cfg[4567] = { 1'b0, 8'h54, 8'h3b}; // CH=0 OP=1
cfg[4568] = { 1'b1, 8'hb8, 8'h5e}; // CH=3 OP=2
cfg[4569] = { 1'b0, 8'h94, 8'he8}; // CH=0 OP=1
cfg[4570] = { 1'b1, 8'h5f, 8'h9a}; // CH=6 OP=3
cfg[4571] = { 1'b0, 8'he7, 8'hf}; // CH=3 OP=1
cfg[4572] = { 1'b1, 8'hea, 8'hf1}; // CH=5 OP=2
cfg[4573] = { 1'b1, 8'h6d, 8'h3e}; // CH=4 OP=3
cfg[4574] = { 1'b0, 8'h5b, 8'hf4}; // CH=3 OP=2
cfg[4575] = { 1'b1, 8'ha1, 8'he9}; // CH=4 OP=0
cfg[4576] = { 1'b1, 8'h6c, 8'h18}; // CH=3 OP=3
cfg[4577] = { 1'b1, 8'ha5, 8'h73}; // CH=4 OP=1
cfg[4578] = { 1'b1, 8'h99, 8'h2c}; // CH=4 OP=2
cfg[4579] = { 1'b0, 8'h34, 8'he7}; // CH=0 OP=1
cfg[4580] = { 1'b1, 8'h7e, 8'h46}; // CH=5 OP=3
cfg[4581] = { 1'b0, 8'h8b, 8'h2d}; // CH=3 OP=2
cfg[4582] = { 1'b1, 8'hb8, 8'h17}; // CH=3 OP=2
cfg[4583] = { 1'b1, 8'ha0, 8'h85}; // CH=3 OP=0
cfg[4584] = { 1'b0, 8'hb0, 8'he0}; // CH=0 OP=0
cfg[4585] = { 1'b1, 8'hf7, 8'h81}; // CH=6 OP=1
cfg[4586] = { 1'b0, 8'h4a, 8'h85}; // CH=2 OP=2
cfg[4587] = { 1'b0, 8'hfc, 8'h2b}; // CH=0 OP=3
cfg[4588] = { 1'b0, 8'h95, 8'h3e}; // CH=1 OP=1
cfg[4589] = { 1'b0, 8'hc9, 8'h25}; // CH=1 OP=2
cfg[4590] = { 1'b1, 8'h48, 8'h6b}; // CH=3 OP=2
cfg[4591] = { 1'b1, 8'hd3, 8'h99}; // CH=6 OP=0
cfg[4592] = { 1'b0, 8'h8c, 8'hb0}; // CH=0 OP=3
cfg[4593] = { 1'b0, 8'h50, 8'h35}; // CH=0 OP=0
cfg[4594] = { 1'b1, 8'h97, 8'hdc}; // CH=6 OP=1
cfg[4595] = { 1'b0, 8'h37, 8'h27}; // CH=3 OP=1
cfg[4596] = { 1'b1, 8'h4b, 8'h71}; // CH=6 OP=2
cfg[4597] = { 1'b0, 8'h8b, 8'h6d}; // CH=3 OP=2
cfg[4598] = { 1'b1, 8'h8b, 8'h3}; // CH=6 OP=2
cfg[4599] = { 1'b0, 8'h4e, 8'hcc}; // CH=2 OP=3
cfg[4600] = { 1'b0, 8'he3, 8'h14}; // CH=3 OP=0
cfg[4601] = { 1'b1, 8'h3c, 8'he8}; // CH=3 OP=3
cfg[4602] = { 1'b1, 8'h96, 8'h74}; // CH=5 OP=1
cfg[4603] = { 1'b1, 8'he6, 8'ha0}; // CH=5 OP=1
cfg[4604] = { 1'b0, 8'ha1, 8'h7d}; // CH=1 OP=0
cfg[4605] = { 1'b1, 8'hd9, 8'h3c}; // CH=4 OP=2
cfg[4606] = { 1'b0, 8'h95, 8'hae}; // CH=1 OP=1
cfg[4607] = { 1'b1, 8'h7a, 8'hb0}; // CH=5 OP=2
cfg[4608] = { 1'b0, 8'h84, 8'h3b}; // CH=0 OP=1
cfg[4609] = { 1'b1, 8'hfa, 8'h8a}; // CH=5 OP=2
cfg[4610] = { 1'b1, 8'he7, 8'h6d}; // CH=6 OP=1
cfg[4611] = { 1'b1, 8'h5b, 8'hc9}; // CH=6 OP=2
cfg[4612] = { 1'b1, 8'hfc, 8'hbe}; // CH=3 OP=3
cfg[4613] = { 1'b1, 8'h79, 8'hc8}; // CH=4 OP=2
cfg[4614] = { 1'b1, 8'hec, 8'h6a}; // CH=3 OP=3
cfg[4615] = { 1'b1, 8'hda, 8'h43}; // CH=5 OP=2
cfg[4616] = { 1'b1, 8'h6f, 8'h67}; // CH=6 OP=3
cfg[4617] = { 1'b1, 8'he9, 8'h17}; // CH=4 OP=2
cfg[4618] = { 1'b1, 8'h6e, 8'h53}; // CH=5 OP=3
cfg[4619] = { 1'b0, 8'h68, 8'hdd}; // CH=0 OP=2
cfg[4620] = { 1'b0, 8'h72, 8'h4a}; // CH=2 OP=0
cfg[4621] = { 1'b1, 8'h3b, 8'hf4}; // CH=6 OP=2
cfg[4622] = { 1'b1, 8'hf9, 8'h33}; // CH=4 OP=2
cfg[4623] = { 1'b1, 8'hc1, 8'h59}; // CH=4 OP=0
cfg[4624] = { 1'b0, 8'hee, 8'h94}; // CH=2 OP=3
cfg[4625] = { 1'b1, 8'hc8, 8'h6e}; // CH=3 OP=2
cfg[4626] = { 1'b1, 8'h38, 8'hd6}; // CH=3 OP=2
cfg[4627] = { 1'b0, 8'hd1, 8'hed}; // CH=1 OP=0
cfg[4628] = { 1'b0, 8'hf8, 8'h8f}; // CH=0 OP=2
cfg[4629] = { 1'b0, 8'h6a, 8'h68}; // CH=2 OP=2
cfg[4630] = { 1'b1, 8'ha5, 8'h5c}; // CH=4 OP=1
cfg[4631] = { 1'b0, 8'h9e, 8'h8f}; // CH=2 OP=3
cfg[4632] = { 1'b1, 8'h5f, 8'he8}; // CH=6 OP=3
cfg[4633] = { 1'b1, 8'h8b, 8'h7c}; // CH=6 OP=2
cfg[4634] = { 1'b1, 8'hf9, 8'h88}; // CH=4 OP=2
cfg[4635] = { 1'b0, 8'hcf, 8'hb9}; // CH=3 OP=3
cfg[4636] = { 1'b0, 8'hbd, 8'h2b}; // CH=1 OP=3
cfg[4637] = { 1'b1, 8'hfd, 8'hfc}; // CH=4 OP=3
cfg[4638] = { 1'b1, 8'h47, 8'h18}; // CH=6 OP=1
cfg[4639] = { 1'b0, 8'hb1, 8'h83}; // CH=1 OP=0
cfg[4640] = { 1'b0, 8'h56, 8'hdf}; // CH=2 OP=1
cfg[4641] = { 1'b0, 8'hf4, 8'h6e}; // CH=0 OP=1
cfg[4642] = { 1'b0, 8'h53, 8'h57}; // CH=3 OP=0
cfg[4643] = { 1'b1, 8'hde, 8'hd3}; // CH=5 OP=3
cfg[4644] = { 1'b1, 8'hd8, 8'h5b}; // CH=3 OP=2
cfg[4645] = { 1'b1, 8'ha7, 8'h14}; // CH=6 OP=1
cfg[4646] = { 1'b1, 8'h64, 8'h3f}; // CH=3 OP=1
cfg[4647] = { 1'b0, 8'h62, 8'h3c}; // CH=2 OP=0
cfg[4648] = { 1'b1, 8'h7d, 8'h54}; // CH=4 OP=3
cfg[4649] = { 1'b0, 8'h3f, 8'hd3}; // CH=3 OP=3
cfg[4650] = { 1'b1, 8'h95, 8'hdf}; // CH=4 OP=1
cfg[4651] = { 1'b1, 8'h89, 8'h4d}; // CH=4 OP=2
cfg[4652] = { 1'b1, 8'hdd, 8'ha4}; // CH=4 OP=3
cfg[4653] = { 1'b1, 8'hbb, 8'h78}; // CH=6 OP=2
cfg[4654] = { 1'b0, 8'h93, 8'hd3}; // CH=3 OP=0
cfg[4655] = { 1'b1, 8'h3b, 8'he8}; // CH=6 OP=2
cfg[4656] = { 1'b0, 8'h9f, 8'h27}; // CH=3 OP=3
cfg[4657] = { 1'b0, 8'hec, 8'h63}; // CH=0 OP=3
cfg[4658] = { 1'b0, 8'h7a, 8'h7e}; // CH=2 OP=2
cfg[4659] = { 1'b1, 8'hba, 8'h7e}; // CH=5 OP=2
cfg[4660] = { 1'b0, 8'h4f, 8'h5d}; // CH=3 OP=3
cfg[4661] = { 1'b1, 8'hd9, 8'hab}; // CH=4 OP=2
cfg[4662] = { 1'b1, 8'hb6, 8'h4f}; // CH=5 OP=1
cfg[4663] = { 1'b0, 8'h71, 8'hc7}; // CH=1 OP=0
cfg[4664] = { 1'b0, 8'h91, 8'h9b}; // CH=1 OP=0
cfg[4665] = { 1'b1, 8'h3d, 8'h40}; // CH=4 OP=3
cfg[4666] = { 1'b0, 8'he1, 8'hdf}; // CH=1 OP=0
cfg[4667] = { 1'b0, 8'hcd, 8'he1}; // CH=1 OP=3
cfg[4668] = { 1'b0, 8'h48, 8'h5f}; // CH=0 OP=2
cfg[4669] = { 1'b1, 8'hc5, 8'hde}; // CH=4 OP=1
cfg[4670] = { 1'b1, 8'h5c, 8'h51}; // CH=3 OP=3
cfg[4671] = { 1'b0, 8'hff, 8'h2a}; // CH=3 OP=3
cfg[4672] = { 1'b0, 8'h45, 8'he0}; // CH=1 OP=1
cfg[4673] = { 1'b1, 8'h63, 8'h52}; // CH=6 OP=0
cfg[4674] = { 1'b0, 8'hf4, 8'h57}; // CH=0 OP=1
cfg[4675] = { 1'b1, 8'h31, 8'h97}; // CH=4 OP=0
cfg[4676] = { 1'b0, 8'hd4, 8'h76}; // CH=0 OP=1
cfg[4677] = { 1'b1, 8'h9a, 8'he0}; // CH=5 OP=2
cfg[4678] = { 1'b1, 8'heb, 8'h28}; // CH=6 OP=2
cfg[4679] = { 1'b1, 8'hb0, 8'h2a}; // CH=3 OP=0
cfg[4680] = { 1'b0, 8'hb7, 8'h7c}; // CH=3 OP=1
cfg[4681] = { 1'b0, 8'hed, 8'hc}; // CH=1 OP=3
cfg[4682] = { 1'b1, 8'hea, 8'h51}; // CH=5 OP=2
cfg[4683] = { 1'b1, 8'h83, 8'hb5}; // CH=6 OP=0
cfg[4684] = { 1'b0, 8'h9e, 8'ha9}; // CH=2 OP=3
cfg[4685] = { 1'b1, 8'h64, 8'hdb}; // CH=3 OP=1
cfg[4686] = { 1'b1, 8'h38, 8'hee}; // CH=3 OP=2
cfg[4687] = { 1'b1, 8'hd2, 8'hce}; // CH=5 OP=0
cfg[4688] = { 1'b0, 8'hbd, 8'hf7}; // CH=1 OP=3
cfg[4689] = { 1'b1, 8'h6d, 8'h21}; // CH=4 OP=3
cfg[4690] = { 1'b1, 8'h7a, 8'h9d}; // CH=5 OP=2
cfg[4691] = { 1'b0, 8'h86, 8'h44}; // CH=2 OP=1
cfg[4692] = { 1'b1, 8'hd7, 8'hcb}; // CH=6 OP=1
cfg[4693] = { 1'b0, 8'h8c, 8'ha4}; // CH=0 OP=3
cfg[4694] = { 1'b1, 8'h36, 8'hd4}; // CH=5 OP=1
cfg[4695] = { 1'b1, 8'hc6, 8'h9b}; // CH=5 OP=1
cfg[4696] = { 1'b0, 8'hfe, 8'hff}; // CH=2 OP=3
cfg[4697] = { 1'b1, 8'hd1, 8'hcd}; // CH=4 OP=0
cfg[4698] = { 1'b1, 8'h8e, 8'hc4}; // CH=5 OP=3
cfg[4699] = { 1'b0, 8'hfc, 8'he6}; // CH=0 OP=3
cfg[4700] = { 1'b0, 8'h76, 8'h83}; // CH=2 OP=1
cfg[4701] = { 1'b0, 8'hfc, 8'hc7}; // CH=0 OP=3
cfg[4702] = { 1'b0, 8'hd3, 8'h92}; // CH=3 OP=0
cfg[4703] = { 1'b0, 8'h60, 8'h36}; // CH=0 OP=0
cfg[4704] = { 1'b1, 8'h96, 8'ha}; // CH=5 OP=1
cfg[4705] = { 1'b0, 8'ha7, 8'ha5}; // CH=3 OP=1
cfg[4706] = { 1'b0, 8'ha6, 8'h7e}; // CH=2 OP=1
cfg[4707] = { 1'b1, 8'h73, 8'heb}; // CH=6 OP=0
cfg[4708] = { 1'b0, 8'h38, 8'ha5}; // CH=0 OP=2
cfg[4709] = { 1'b0, 8'h8e, 8'h3f}; // CH=2 OP=3
cfg[4710] = { 1'b1, 8'h40, 8'ha1}; // CH=3 OP=0
cfg[4711] = { 1'b1, 8'h4a, 8'h0}; // CH=5 OP=2
cfg[4712] = { 1'b1, 8'h94, 8'hd4}; // CH=3 OP=1
cfg[4713] = { 1'b0, 8'ha1, 8'h34}; // CH=1 OP=0
cfg[4714] = { 1'b0, 8'he2, 8'hca}; // CH=2 OP=0
cfg[4715] = { 1'b1, 8'h60, 8'h44}; // CH=3 OP=0
cfg[4716] = { 1'b1, 8'h4b, 8'h77}; // CH=6 OP=2
cfg[4717] = { 1'b0, 8'hf0, 8'h7b}; // CH=0 OP=0
cfg[4718] = { 1'b0, 8'h30, 8'hd}; // CH=0 OP=0
cfg[4719] = { 1'b0, 8'hbb, 8'h9c}; // CH=3 OP=2
cfg[4720] = { 1'b0, 8'hfb, 8'ha0}; // CH=3 OP=2
cfg[4721] = { 1'b1, 8'h45, 8'ha1}; // CH=4 OP=1
cfg[4722] = { 1'b0, 8'hd9, 8'h75}; // CH=1 OP=2
cfg[4723] = { 1'b0, 8'h7a, 8'ha9}; // CH=2 OP=2
cfg[4724] = { 1'b1, 8'h8a, 8'h73}; // CH=5 OP=2
cfg[4725] = { 1'b1, 8'hce, 8'he4}; // CH=5 OP=3
cfg[4726] = { 1'b1, 8'h45, 8'hfb}; // CH=4 OP=1
cfg[4727] = { 1'b0, 8'hc0, 8'h85}; // CH=0 OP=0
cfg[4728] = { 1'b1, 8'hcd, 8'h48}; // CH=4 OP=3
cfg[4729] = { 1'b1, 8'h69, 8'h28}; // CH=4 OP=2
cfg[4730] = { 1'b0, 8'hba, 8'haa}; // CH=2 OP=2
cfg[4731] = { 1'b1, 8'hff, 8'hab}; // CH=6 OP=3
cfg[4732] = { 1'b0, 8'hd9, 8'h20}; // CH=1 OP=2
cfg[4733] = { 1'b0, 8'h53, 8'hc9}; // CH=3 OP=0
cfg[4734] = { 1'b1, 8'hdd, 8'h3c}; // CH=4 OP=3
cfg[4735] = { 1'b0, 8'hab, 8'h20}; // CH=3 OP=2
cfg[4736] = { 1'b1, 8'hf0, 8'h1b}; // CH=3 OP=0
cfg[4737] = { 1'b0, 8'hb0, 8'ha0}; // CH=0 OP=0
cfg[4738] = { 1'b1, 8'h7e, 8'he8}; // CH=5 OP=3
cfg[4739] = { 1'b0, 8'he7, 8'h11}; // CH=3 OP=1
cfg[4740] = { 1'b0, 8'hf1, 8'hbb}; // CH=1 OP=0
cfg[4741] = { 1'b0, 8'h9c, 8'h51}; // CH=0 OP=3
cfg[4742] = { 1'b0, 8'hbc, 8'hcd}; // CH=0 OP=3
cfg[4743] = { 1'b1, 8'h85, 8'h61}; // CH=4 OP=1
cfg[4744] = { 1'b0, 8'hc1, 8'h4b}; // CH=1 OP=0
cfg[4745] = { 1'b0, 8'he1, 8'h6b}; // CH=1 OP=0
cfg[4746] = { 1'b1, 8'hfc, 8'h23}; // CH=3 OP=3
cfg[4747] = { 1'b0, 8'h9d, 8'hbd}; // CH=1 OP=3
cfg[4748] = { 1'b0, 8'h85, 8'h2a}; // CH=1 OP=1
cfg[4749] = { 1'b0, 8'h96, 8'h9a}; // CH=2 OP=1
cfg[4750] = { 1'b0, 8'h52, 8'hc8}; // CH=2 OP=0
cfg[4751] = { 1'b1, 8'ha3, 8'hb1}; // CH=6 OP=0
cfg[4752] = { 1'b0, 8'h70, 8'h99}; // CH=0 OP=0
cfg[4753] = { 1'b0, 8'hd1, 8'h5a}; // CH=1 OP=0
cfg[4754] = { 1'b0, 8'h35, 8'h6e}; // CH=1 OP=1
cfg[4755] = { 1'b0, 8'hfe, 8'h88}; // CH=2 OP=3
cfg[4756] = { 1'b1, 8'h8c, 8'h13}; // CH=3 OP=3
cfg[4757] = { 1'b0, 8'hca, 8'hb0}; // CH=2 OP=2
cfg[4758] = { 1'b0, 8'h87, 8'h36}; // CH=3 OP=1
cfg[4759] = { 1'b0, 8'hf4, 8'hcc}; // CH=0 OP=1
cfg[4760] = { 1'b0, 8'ha5, 8'hc0}; // CH=1 OP=1
cfg[4761] = { 1'b1, 8'h3e, 8'hf2}; // CH=5 OP=3
cfg[4762] = { 1'b1, 8'h98, 8'he1}; // CH=3 OP=2
cfg[4763] = { 1'b1, 8'h8a, 8'h55}; // CH=5 OP=2
cfg[4764] = { 1'b1, 8'ha1, 8'ha7}; // CH=4 OP=0
cfg[4765] = { 1'b1, 8'hb5, 8'h52}; // CH=4 OP=1
cfg[4766] = { 1'b1, 8'h65, 8'hba}; // CH=4 OP=1
cfg[4767] = { 1'b0, 8'h9b, 8'h4c}; // CH=3 OP=2
cfg[4768] = { 1'b1, 8'h68, 8'h78}; // CH=3 OP=2
cfg[4769] = { 1'b0, 8'h86, 8'h6d}; // CH=2 OP=1
cfg[4770] = { 1'b0, 8'h48, 8'h12}; // CH=0 OP=2
cfg[4771] = { 1'b1, 8'h79, 8'h51}; // CH=4 OP=2
cfg[4772] = { 1'b0, 8'h7c, 8'he9}; // CH=0 OP=3
cfg[4773] = { 1'b1, 8'h9c, 8'hf0}; // CH=3 OP=3
cfg[4774] = { 1'b1, 8'h43, 8'h58}; // CH=6 OP=0
cfg[4775] = { 1'b1, 8'h96, 8'hbd}; // CH=5 OP=1
cfg[4776] = { 1'b0, 8'h50, 8'haf}; // CH=0 OP=0
cfg[4777] = { 1'b1, 8'h9d, 8'h6b}; // CH=4 OP=3
cfg[4778] = { 1'b1, 8'ha1, 8'hae}; // CH=4 OP=0
cfg[4779] = { 1'b0, 8'h4a, 8'h82}; // CH=2 OP=2
cfg[4780] = { 1'b1, 8'h6b, 8'h6f}; // CH=6 OP=2
cfg[4781] = { 1'b0, 8'h6d, 8'he9}; // CH=1 OP=3
cfg[4782] = { 1'b1, 8'hc4, 8'h65}; // CH=3 OP=1
cfg[4783] = { 1'b0, 8'ha6, 8'h1}; // CH=2 OP=1
cfg[4784] = { 1'b0, 8'hd5, 8'h45}; // CH=1 OP=1
cfg[4785] = { 1'b1, 8'h84, 8'h61}; // CH=3 OP=1
cfg[4786] = { 1'b1, 8'hef, 8'hfe}; // CH=6 OP=3
cfg[4787] = { 1'b0, 8'h9d, 8'h37}; // CH=1 OP=3
cfg[4788] = { 1'b0, 8'hb9, 8'hd8}; // CH=1 OP=2
cfg[4789] = { 1'b0, 8'hf5, 8'h0}; // CH=1 OP=1
cfg[4790] = { 1'b1, 8'hdb, 8'h6f}; // CH=6 OP=2
cfg[4791] = { 1'b0, 8'hab, 8'hdd}; // CH=3 OP=2
cfg[4792] = { 1'b0, 8'h6b, 8'ha1}; // CH=3 OP=2
cfg[4793] = { 1'b1, 8'h83, 8'h47}; // CH=6 OP=0
cfg[4794] = { 1'b0, 8'h58, 8'h70}; // CH=0 OP=2
cfg[4795] = { 1'b1, 8'hdd, 8'hd1}; // CH=4 OP=3
cfg[4796] = { 1'b1, 8'hcc, 8'hd0}; // CH=3 OP=3
cfg[4797] = { 1'b1, 8'h6a, 8'h7}; // CH=5 OP=2
cfg[4798] = { 1'b1, 8'he0, 8'he0}; // CH=3 OP=0
cfg[4799] = { 1'b1, 8'h4f, 8'h7}; // CH=6 OP=3
cfg[4800] = { 1'b1, 8'ha8, 8'he3}; // CH=3 OP=2
cfg[4801] = { 1'b0, 8'h66, 8'h8e}; // CH=2 OP=1
cfg[4802] = { 1'b1, 8'h5d, 8'hf9}; // CH=4 OP=3
cfg[4803] = { 1'b0, 8'hcd, 8'h2a}; // CH=1 OP=3
cfg[4804] = { 1'b0, 8'h9f, 8'h9}; // CH=3 OP=3
cfg[4805] = { 1'b1, 8'h6f, 8'h14}; // CH=6 OP=3
cfg[4806] = { 1'b0, 8'h76, 8'he8}; // CH=2 OP=1
cfg[4807] = { 1'b0, 8'h56, 8'h99}; // CH=2 OP=1
cfg[4808] = { 1'b1, 8'h36, 8'hab}; // CH=5 OP=1
cfg[4809] = { 1'b1, 8'h86, 8'hb3}; // CH=5 OP=1
cfg[4810] = { 1'b0, 8'h3e, 8'h96}; // CH=2 OP=3
cfg[4811] = { 1'b0, 8'h53, 8'h94}; // CH=3 OP=0
cfg[4812] = { 1'b1, 8'hb0, 8'hb9}; // CH=3 OP=0
cfg[4813] = { 1'b1, 8'h7e, 8'he3}; // CH=5 OP=3
cfg[4814] = { 1'b1, 8'h8c, 8'hed}; // CH=3 OP=3
cfg[4815] = { 1'b1, 8'h85, 8'he9}; // CH=4 OP=1
cfg[4816] = { 1'b1, 8'h90, 8'h59}; // CH=3 OP=0
cfg[4817] = { 1'b0, 8'hc3, 8'h8f}; // CH=3 OP=0
cfg[4818] = { 1'b1, 8'h8d, 8'h15}; // CH=4 OP=3
cfg[4819] = { 1'b1, 8'hcb, 8'h43}; // CH=6 OP=2
cfg[4820] = { 1'b1, 8'hb8, 8'hd7}; // CH=3 OP=2
cfg[4821] = { 1'b1, 8'h51, 8'hcf}; // CH=4 OP=0
cfg[4822] = { 1'b0, 8'hbf, 8'h4d}; // CH=3 OP=3
cfg[4823] = { 1'b1, 8'hde, 8'h6a}; // CH=5 OP=3
cfg[4824] = { 1'b1, 8'h7b, 8'hf6}; // CH=6 OP=2
cfg[4825] = { 1'b0, 8'hcf, 8'hf9}; // CH=3 OP=3
cfg[4826] = { 1'b0, 8'hfe, 8'h90}; // CH=2 OP=3
cfg[4827] = { 1'b1, 8'hdf, 8'h54}; // CH=6 OP=3
cfg[4828] = { 1'b1, 8'h57, 8'he1}; // CH=6 OP=1
cfg[4829] = { 1'b0, 8'hf2, 8'had}; // CH=2 OP=0
cfg[4830] = { 1'b0, 8'hab, 8'hcc}; // CH=3 OP=2
cfg[4831] = { 1'b1, 8'hfc, 8'h9b}; // CH=3 OP=3
cfg[4832] = { 1'b1, 8'hbb, 8'he9}; // CH=6 OP=2
cfg[4833] = { 1'b1, 8'h99, 8'h53}; // CH=4 OP=2
cfg[4834] = { 1'b0, 8'h43, 8'h4a}; // CH=3 OP=0
cfg[4835] = { 1'b0, 8'h95, 8'hf8}; // CH=1 OP=1
cfg[4836] = { 1'b1, 8'h76, 8'hf6}; // CH=5 OP=1
cfg[4837] = { 1'b1, 8'h6d, 8'hd5}; // CH=4 OP=3
cfg[4838] = { 1'b0, 8'ha8, 8'h2c}; // CH=0 OP=2
cfg[4839] = { 1'b1, 8'hba, 8'h1f}; // CH=5 OP=2
cfg[4840] = { 1'b1, 8'h5d, 8'hca}; // CH=4 OP=3
cfg[4841] = { 1'b1, 8'h74, 8'hc6}; // CH=3 OP=1
cfg[4842] = { 1'b0, 8'hed, 8'h82}; // CH=1 OP=3
cfg[4843] = { 1'b1, 8'hc9, 8'h1b}; // CH=4 OP=2
cfg[4844] = { 1'b1, 8'hf2, 8'h30}; // CH=5 OP=0
cfg[4845] = { 1'b0, 8'hea, 8'h44}; // CH=2 OP=2
cfg[4846] = { 1'b1, 8'he0, 8'he9}; // CH=3 OP=0
cfg[4847] = { 1'b0, 8'hb5, 8'he2}; // CH=1 OP=1
cfg[4848] = { 1'b1, 8'he2, 8'hbd}; // CH=5 OP=0
cfg[4849] = { 1'b1, 8'h93, 8'h44}; // CH=6 OP=0
cfg[4850] = { 1'b0, 8'hf0, 8'hcb}; // CH=0 OP=0
cfg[4851] = { 1'b1, 8'h65, 8'h91}; // CH=4 OP=1
cfg[4852] = { 1'b1, 8'h52, 8'h13}; // CH=5 OP=0
cfg[4853] = { 1'b0, 8'h5f, 8'h2f}; // CH=3 OP=3
cfg[4854] = { 1'b0, 8'ha3, 8'hb8}; // CH=3 OP=0
cfg[4855] = { 1'b0, 8'h8d, 8'h6}; // CH=1 OP=3
cfg[4856] = { 1'b0, 8'h6f, 8'hca}; // CH=3 OP=3
cfg[4857] = { 1'b1, 8'h6f, 8'hfb}; // CH=6 OP=3
cfg[4858] = { 1'b1, 8'h70, 8'h71}; // CH=3 OP=0
cfg[4859] = { 1'b0, 8'h3b, 8'h9}; // CH=3 OP=2
cfg[4860] = { 1'b1, 8'hcd, 8'h90}; // CH=4 OP=3
cfg[4861] = { 1'b0, 8'he0, 8'hef}; // CH=0 OP=0
cfg[4862] = { 1'b0, 8'h79, 8'h79}; // CH=1 OP=2
cfg[4863] = { 1'b0, 8'h32, 8'h3a}; // CH=2 OP=0
cfg[4864] = { 1'b0, 8'h38, 8'h32}; // CH=0 OP=2
cfg[4865] = { 1'b1, 8'h98, 8'ha}; // CH=3 OP=2
cfg[4866] = { 1'b1, 8'hd2, 8'h3b}; // CH=5 OP=0
cfg[4867] = { 1'b0, 8'h3b, 8'h78}; // CH=3 OP=2
cfg[4868] = { 1'b1, 8'h94, 8'hb3}; // CH=3 OP=1
cfg[4869] = { 1'b1, 8'h52, 8'h80}; // CH=5 OP=0
cfg[4870] = { 1'b0, 8'h62, 8'h61}; // CH=2 OP=0
cfg[4871] = { 1'b1, 8'h8f, 8'h70}; // CH=6 OP=3
cfg[4872] = { 1'b1, 8'hc9, 8'hdf}; // CH=4 OP=2
cfg[4873] = { 1'b1, 8'hfc, 8'hf1}; // CH=3 OP=3
cfg[4874] = { 1'b1, 8'h93, 8'h90}; // CH=6 OP=0
cfg[4875] = { 1'b0, 8'h90, 8'h9e}; // CH=0 OP=0
cfg[4876] = { 1'b1, 8'h63, 8'ha6}; // CH=6 OP=0
cfg[4877] = { 1'b1, 8'h9e, 8'h1e}; // CH=5 OP=3
cfg[4878] = { 1'b0, 8'h32, 8'hd1}; // CH=2 OP=0
cfg[4879] = { 1'b1, 8'h84, 8'h52}; // CH=3 OP=1
cfg[4880] = { 1'b1, 8'he6, 8'hb3}; // CH=5 OP=1
cfg[4881] = { 1'b1, 8'h75, 8'h23}; // CH=4 OP=1
cfg[4882] = { 1'b0, 8'h3f, 8'h2}; // CH=3 OP=3
cfg[4883] = { 1'b1, 8'h3b, 8'hf3}; // CH=6 OP=2
cfg[4884] = { 1'b0, 8'h41, 8'h83}; // CH=1 OP=0
cfg[4885] = { 1'b1, 8'he0, 8'h22}; // CH=3 OP=0
cfg[4886] = { 1'b1, 8'h86, 8'hfb}; // CH=5 OP=1
cfg[4887] = { 1'b0, 8'ha4, 8'h81}; // CH=0 OP=1
cfg[4888] = { 1'b0, 8'h75, 8'hbb}; // CH=1 OP=1
cfg[4889] = { 1'b0, 8'hc7, 8'h3b}; // CH=3 OP=1
cfg[4890] = { 1'b0, 8'h7a, 8'hee}; // CH=2 OP=2
cfg[4891] = { 1'b1, 8'h9e, 8'h4f}; // CH=5 OP=3
cfg[4892] = { 1'b0, 8'ha0, 8'hd7}; // CH=0 OP=0
cfg[4893] = { 1'b1, 8'h94, 8'hb8}; // CH=3 OP=1
cfg[4894] = { 1'b0, 8'h64, 8'h2a}; // CH=0 OP=1
cfg[4895] = { 1'b1, 8'h44, 8'h39}; // CH=3 OP=1
cfg[4896] = { 1'b1, 8'hca, 8'h35}; // CH=5 OP=2
cfg[4897] = { 1'b1, 8'h6e, 8'hb6}; // CH=5 OP=3
cfg[4898] = { 1'b0, 8'he3, 8'h71}; // CH=3 OP=0
cfg[4899] = { 1'b0, 8'hab, 8'hac}; // CH=3 OP=2
cfg[4900] = { 1'b1, 8'h9c, 8'h9b}; // CH=3 OP=3
cfg[4901] = { 1'b0, 8'h44, 8'hc3}; // CH=0 OP=1
cfg[4902] = { 1'b0, 8'h7a, 8'h64}; // CH=2 OP=2
cfg[4903] = { 1'b0, 8'ha5, 8'h4e}; // CH=1 OP=1
cfg[4904] = { 1'b1, 8'hd4, 8'hb2}; // CH=3 OP=1
cfg[4905] = { 1'b1, 8'h99, 8'hf6}; // CH=4 OP=2
cfg[4906] = { 1'b0, 8'h57, 8'hc0}; // CH=3 OP=1
cfg[4907] = { 1'b0, 8'hab, 8'h2e}; // CH=3 OP=2
cfg[4908] = { 1'b1, 8'hc7, 8'h12}; // CH=6 OP=1
cfg[4909] = { 1'b0, 8'h30, 8'hbd}; // CH=0 OP=0
cfg[4910] = { 1'b1, 8'hcc, 8'he2}; // CH=3 OP=3
cfg[4911] = { 1'b1, 8'h99, 8'ha6}; // CH=4 OP=2
cfg[4912] = { 1'b0, 8'h8b, 8'h3d}; // CH=3 OP=2
cfg[4913] = { 1'b1, 8'h3e, 8'h11}; // CH=5 OP=3
cfg[4914] = { 1'b1, 8'h34, 8'h5a}; // CH=3 OP=1
cfg[4915] = { 1'b1, 8'hf5, 8'hd8}; // CH=4 OP=1
cfg[4916] = { 1'b0, 8'hb2, 8'hc}; // CH=2 OP=0
cfg[4917] = { 1'b1, 8'hf2, 8'hf0}; // CH=5 OP=0
cfg[4918] = { 1'b1, 8'hd5, 8'hf1}; // CH=4 OP=1
cfg[4919] = { 1'b1, 8'h7b, 8'hc8}; // CH=6 OP=2
cfg[4920] = { 1'b0, 8'h85, 8'h62}; // CH=1 OP=1
cfg[4921] = { 1'b1, 8'h87, 8'h76}; // CH=6 OP=1
cfg[4922] = { 1'b1, 8'h98, 8'h2f}; // CH=3 OP=2
cfg[4923] = { 1'b1, 8'hf3, 8'hbc}; // CH=6 OP=0
cfg[4924] = { 1'b1, 8'hcb, 8'he3}; // CH=6 OP=2
cfg[4925] = { 1'b0, 8'hd8, 8'h61}; // CH=0 OP=2
cfg[4926] = { 1'b0, 8'h8a, 8'h8a}; // CH=2 OP=2
cfg[4927] = { 1'b1, 8'h8e, 8'h7b}; // CH=5 OP=3
cfg[4928] = { 1'b0, 8'h7f, 8'h9c}; // CH=3 OP=3
cfg[4929] = { 1'b1, 8'h47, 8'h89}; // CH=6 OP=1
cfg[4930] = { 1'b0, 8'ha9, 8'h88}; // CH=1 OP=2
cfg[4931] = { 1'b1, 8'hd6, 8'hc3}; // CH=5 OP=1
cfg[4932] = { 1'b0, 8'h6e, 8'h4e}; // CH=2 OP=3
cfg[4933] = { 1'b1, 8'h61, 8'hb}; // CH=4 OP=0
cfg[4934] = { 1'b1, 8'hf7, 8'hee}; // CH=6 OP=1
cfg[4935] = { 1'b0, 8'h49, 8'h5}; // CH=1 OP=2
cfg[4936] = { 1'b0, 8'hd1, 8'h8f}; // CH=1 OP=0
cfg[4937] = { 1'b1, 8'h4b, 8'h1d}; // CH=6 OP=2
cfg[4938] = { 1'b1, 8'h9a, 8'h9c}; // CH=5 OP=2
cfg[4939] = { 1'b1, 8'h64, 8'he3}; // CH=3 OP=1
cfg[4940] = { 1'b1, 8'hb3, 8'h8d}; // CH=6 OP=0
cfg[4941] = { 1'b0, 8'h89, 8'hac}; // CH=1 OP=2
cfg[4942] = { 1'b1, 8'hf7, 8'hfb}; // CH=6 OP=1
cfg[4943] = { 1'b0, 8'h59, 8'h6}; // CH=1 OP=2
cfg[4944] = { 1'b1, 8'h86, 8'hf4}; // CH=5 OP=1
cfg[4945] = { 1'b1, 8'h8b, 8'h44}; // CH=6 OP=2
cfg[4946] = { 1'b0, 8'hbb, 8'h1f}; // CH=3 OP=2
cfg[4947] = { 1'b0, 8'h66, 8'h37}; // CH=2 OP=1
cfg[4948] = { 1'b1, 8'he1, 8'ha0}; // CH=4 OP=0
cfg[4949] = { 1'b0, 8'he4, 8'h4}; // CH=0 OP=1
cfg[4950] = { 1'b1, 8'haa, 8'hb7}; // CH=5 OP=2
cfg[4951] = { 1'b0, 8'hfb, 8'h40}; // CH=3 OP=2
cfg[4952] = { 1'b1, 8'hdc, 8'h38}; // CH=3 OP=3
cfg[4953] = { 1'b1, 8'h85, 8'h91}; // CH=4 OP=1
cfg[4954] = { 1'b1, 8'ha2, 8'h17}; // CH=5 OP=0
cfg[4955] = { 1'b1, 8'hbc, 8'h49}; // CH=3 OP=3
cfg[4956] = { 1'b0, 8'hf3, 8'hbd}; // CH=3 OP=0
cfg[4957] = { 1'b1, 8'hc6, 8'h23}; // CH=5 OP=1
cfg[4958] = { 1'b1, 8'h7c, 8'h4}; // CH=3 OP=3
cfg[4959] = { 1'b0, 8'hc0, 8'he8}; // CH=0 OP=0
cfg[4960] = { 1'b1, 8'hb0, 8'h93}; // CH=3 OP=0
cfg[4961] = { 1'b0, 8'h9b, 8'h8e}; // CH=3 OP=2
cfg[4962] = { 1'b0, 8'h8c, 8'h6a}; // CH=0 OP=3
cfg[4963] = { 1'b1, 8'h71, 8'hf0}; // CH=4 OP=0
cfg[4964] = { 1'b0, 8'h9b, 8'h16}; // CH=3 OP=2
cfg[4965] = { 1'b0, 8'he4, 8'h27}; // CH=0 OP=1
cfg[4966] = { 1'b0, 8'ha2, 8'hf4}; // CH=2 OP=0
cfg[4967] = { 1'b1, 8'hc5, 8'hc7}; // CH=4 OP=1
cfg[4968] = { 1'b1, 8'hca, 8'h3a}; // CH=5 OP=2
cfg[4969] = { 1'b1, 8'hb2, 8'hb2}; // CH=5 OP=0
cfg[4970] = { 1'b1, 8'h45, 8'he2}; // CH=4 OP=1
cfg[4971] = { 1'b1, 8'hd4, 8'h52}; // CH=3 OP=1
cfg[4972] = { 1'b0, 8'h3e, 8'hfa}; // CH=2 OP=3
cfg[4973] = { 1'b0, 8'hec, 8'h33}; // CH=0 OP=3
cfg[4974] = { 1'b1, 8'h87, 8'h45}; // CH=6 OP=1
cfg[4975] = { 1'b1, 8'h6c, 8'h6c}; // CH=3 OP=3
cfg[4976] = { 1'b1, 8'hc4, 8'h60}; // CH=3 OP=1
cfg[4977] = { 1'b1, 8'h62, 8'hd3}; // CH=5 OP=0
cfg[4978] = { 1'b1, 8'h50, 8'he}; // CH=3 OP=0
cfg[4979] = { 1'b0, 8'h95, 8'hf6}; // CH=1 OP=1
cfg[4980] = { 1'b1, 8'h69, 8'h48}; // CH=4 OP=2
cfg[4981] = { 1'b0, 8'ha8, 8'h42}; // CH=0 OP=2
cfg[4982] = { 1'b0, 8'hd6, 8'h75}; // CH=2 OP=1
cfg[4983] = { 1'b0, 8'he2, 8'hf8}; // CH=2 OP=0
cfg[4984] = { 1'b1, 8'h4e, 8'h88}; // CH=5 OP=3
cfg[4985] = { 1'b0, 8'h5c, 8'he8}; // CH=0 OP=3
cfg[4986] = { 1'b0, 8'h7f, 8'h10}; // CH=3 OP=3
cfg[4987] = { 1'b0, 8'h8e, 8'hcd}; // CH=2 OP=3
cfg[4988] = { 1'b0, 8'h40, 8'h1d}; // CH=0 OP=0
cfg[4989] = { 1'b1, 8'h45, 8'hb2}; // CH=4 OP=1
cfg[4990] = { 1'b1, 8'h39, 8'h1c}; // CH=4 OP=2
cfg[4991] = { 1'b0, 8'ha8, 8'hc4}; // CH=0 OP=2
cfg[4992] = { 1'b1, 8'h76, 8'h9a}; // CH=5 OP=1
cfg[4993] = { 1'b0, 8'he3, 8'he4}; // CH=3 OP=0
cfg[4994] = { 1'b0, 8'h74, 8'h32}; // CH=0 OP=1
cfg[4995] = { 1'b0, 8'hc8, 8'h8e}; // CH=0 OP=2
cfg[4996] = { 1'b0, 8'h48, 8'hbe}; // CH=0 OP=2
cfg[4997] = { 1'b0, 8'hd6, 8'h8b}; // CH=2 OP=1
cfg[4998] = { 1'b1, 8'hac, 8'ha8}; // CH=3 OP=3
cfg[4999] = { 1'b0, 8'h71, 8'h5b}; // CH=1 OP=0

cfg[5000] = { 1'b0, 8'h0, 8'h00 }; // done
