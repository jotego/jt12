cfg[0] = { 1'b0, 8'ha4, 8'h0}; // CH=0 OP=1
cfg[1] = { 1'b0, 8'h30, 8'h67}; // CH=0 OP=0
cfg[2] = { 1'b0, 8'h31, 8'hc6}; // CH=1 OP=0
cfg[3] = { 1'b0, 8'h32, 8'h69}; // CH=2 OP=0
cfg[4] = { 1'b1, 8'h30, 8'h73}; // CH=3 OP=0
cfg[5] = { 1'b1, 8'h31, 8'h51}; // CH=4 OP=0
cfg[6] = { 1'b1, 8'h32, 8'hff}; // CH=5 OP=0
cfg[7] = { 1'b0, 8'h34, 8'h4a}; // CH=0 OP=1
cfg[8] = { 1'b0, 8'h35, 8'hec}; // CH=1 OP=1
cfg[9] = { 1'b0, 8'h36, 8'h29}; // CH=2 OP=1
cfg[10] = { 1'b1, 8'h34, 8'hcd}; // CH=3 OP=1
cfg[11] = { 1'b1, 8'h35, 8'hba}; // CH=4 OP=1
cfg[12] = { 1'b1, 8'h36, 8'hab}; // CH=5 OP=1
cfg[13] = { 1'b0, 8'h38, 8'hf2}; // CH=0 OP=2
cfg[14] = { 1'b0, 8'h39, 8'hfb}; // CH=1 OP=2
cfg[15] = { 1'b0, 8'h3a, 8'he3}; // CH=2 OP=2
cfg[16] = { 1'b1, 8'h38, 8'h46}; // CH=3 OP=2
cfg[17] = { 1'b1, 8'h39, 8'h7c}; // CH=4 OP=2
cfg[18] = { 1'b1, 8'h3a, 8'hc2}; // CH=5 OP=2
cfg[19] = { 1'b0, 8'h3c, 8'h54}; // CH=0 OP=3
cfg[20] = { 1'b0, 8'h3d, 8'hf8}; // CH=1 OP=3
cfg[21] = { 1'b0, 8'h3e, 8'h1b}; // CH=2 OP=3
cfg[22] = { 1'b1, 8'h3c, 8'he8}; // CH=3 OP=3
cfg[23] = { 1'b1, 8'h3d, 8'he7}; // CH=4 OP=3
cfg[24] = { 1'b1, 8'h3e, 8'h8d}; // CH=5 OP=3
cfg[25] = { 1'b0, 8'h40, 8'h76}; // CH=0 OP=0
cfg[26] = { 1'b0, 8'h41, 8'h5a}; // CH=1 OP=0
cfg[27] = { 1'b0, 8'h42, 8'h2e}; // CH=2 OP=0
cfg[28] = { 1'b1, 8'h40, 8'h63}; // CH=3 OP=0
cfg[29] = { 1'b1, 8'h41, 8'h33}; // CH=4 OP=0
cfg[30] = { 1'b1, 8'h42, 8'h9f}; // CH=5 OP=0
cfg[31] = { 1'b0, 8'h44, 8'hc9}; // CH=0 OP=1
cfg[32] = { 1'b0, 8'h45, 8'h9a}; // CH=1 OP=1
cfg[33] = { 1'b0, 8'h46, 8'h66}; // CH=2 OP=1
cfg[34] = { 1'b1, 8'h44, 8'h32}; // CH=3 OP=1
cfg[35] = { 1'b1, 8'h45, 8'hd}; // CH=4 OP=1
cfg[36] = { 1'b1, 8'h46, 8'hb7}; // CH=5 OP=1
cfg[37] = { 1'b0, 8'h48, 8'h31}; // CH=0 OP=2
cfg[38] = { 1'b0, 8'h49, 8'h58}; // CH=1 OP=2
cfg[39] = { 1'b0, 8'h4a, 8'ha3}; // CH=2 OP=2
cfg[40] = { 1'b1, 8'h48, 8'h5a}; // CH=3 OP=2
cfg[41] = { 1'b1, 8'h49, 8'h25}; // CH=4 OP=2
cfg[42] = { 1'b1, 8'h4a, 8'h5d}; // CH=5 OP=2
cfg[43] = { 1'b0, 8'h4c, 8'h5}; // CH=0 OP=3
cfg[44] = { 1'b0, 8'h4d, 8'h17}; // CH=1 OP=3
cfg[45] = { 1'b0, 8'h4e, 8'h58}; // CH=2 OP=3
cfg[46] = { 1'b1, 8'h4c, 8'he9}; // CH=3 OP=3
cfg[47] = { 1'b1, 8'h4d, 8'h5e}; // CH=4 OP=3
cfg[48] = { 1'b1, 8'h4e, 8'hd4}; // CH=5 OP=3
cfg[49] = { 1'b0, 8'h50, 8'hab}; // CH=0 OP=0
cfg[50] = { 1'b0, 8'h51, 8'hb2}; // CH=1 OP=0
cfg[51] = { 1'b0, 8'h52, 8'hcd}; // CH=2 OP=0
cfg[52] = { 1'b1, 8'h50, 8'hc6}; // CH=3 OP=0
cfg[53] = { 1'b1, 8'h51, 8'h9b}; // CH=4 OP=0
cfg[54] = { 1'b1, 8'h52, 8'hb4}; // CH=5 OP=0
cfg[55] = { 1'b0, 8'h54, 8'h54}; // CH=0 OP=1
cfg[56] = { 1'b0, 8'h55, 8'h11}; // CH=1 OP=1
cfg[57] = { 1'b0, 8'h56, 8'he}; // CH=2 OP=1
cfg[58] = { 1'b1, 8'h54, 8'h82}; // CH=3 OP=1
cfg[59] = { 1'b1, 8'h55, 8'h74}; // CH=4 OP=1
cfg[60] = { 1'b1, 8'h56, 8'h41}; // CH=5 OP=1
cfg[61] = { 1'b0, 8'h58, 8'h21}; // CH=0 OP=2
cfg[62] = { 1'b0, 8'h59, 8'h3d}; // CH=1 OP=2
cfg[63] = { 1'b0, 8'h5a, 8'hdc}; // CH=2 OP=2
cfg[64] = { 1'b1, 8'h58, 8'h87}; // CH=3 OP=2
cfg[65] = { 1'b1, 8'h59, 8'h70}; // CH=4 OP=2
cfg[66] = { 1'b1, 8'h5a, 8'he9}; // CH=5 OP=2
cfg[67] = { 1'b0, 8'h5c, 8'h3e}; // CH=0 OP=3
cfg[68] = { 1'b0, 8'h5d, 8'ha1}; // CH=1 OP=3
cfg[69] = { 1'b0, 8'h5e, 8'h41}; // CH=2 OP=3
cfg[70] = { 1'b1, 8'h5c, 8'he1}; // CH=3 OP=3
cfg[71] = { 1'b1, 8'h5d, 8'hfc}; // CH=4 OP=3
cfg[72] = { 1'b1, 8'h5e, 8'h67}; // CH=5 OP=3
cfg[73] = { 1'b0, 8'h60, 8'h3e}; // CH=0 OP=0
cfg[74] = { 1'b0, 8'h61, 8'h1}; // CH=1 OP=0
cfg[75] = { 1'b0, 8'h62, 8'h7e}; // CH=2 OP=0
cfg[76] = { 1'b1, 8'h60, 8'h97}; // CH=3 OP=0
cfg[77] = { 1'b1, 8'h61, 8'hea}; // CH=4 OP=0
cfg[78] = { 1'b1, 8'h62, 8'hdc}; // CH=5 OP=0
cfg[79] = { 1'b0, 8'h64, 8'h6b}; // CH=0 OP=1
cfg[80] = { 1'b0, 8'h65, 8'h96}; // CH=1 OP=1
cfg[81] = { 1'b0, 8'h66, 8'h8f}; // CH=2 OP=1
cfg[82] = { 1'b1, 8'h64, 8'h38}; // CH=3 OP=1
cfg[83] = { 1'b1, 8'h65, 8'h5c}; // CH=4 OP=1
cfg[84] = { 1'b1, 8'h66, 8'h2a}; // CH=5 OP=1
cfg[85] = { 1'b0, 8'h68, 8'hec}; // CH=0 OP=2
cfg[86] = { 1'b0, 8'h69, 8'hb0}; // CH=1 OP=2
cfg[87] = { 1'b0, 8'h6a, 8'h3b}; // CH=2 OP=2
cfg[88] = { 1'b1, 8'h68, 8'hfb}; // CH=3 OP=2
cfg[89] = { 1'b1, 8'h69, 8'h32}; // CH=4 OP=2
cfg[90] = { 1'b1, 8'h6a, 8'haf}; // CH=5 OP=2
cfg[91] = { 1'b0, 8'h6c, 8'h3c}; // CH=0 OP=3
cfg[92] = { 1'b0, 8'h6d, 8'h54}; // CH=1 OP=3
cfg[93] = { 1'b0, 8'h6e, 8'hec}; // CH=2 OP=3
cfg[94] = { 1'b1, 8'h6c, 8'h18}; // CH=3 OP=3
cfg[95] = { 1'b1, 8'h6d, 8'hdb}; // CH=4 OP=3
cfg[96] = { 1'b1, 8'h6e, 8'h5c}; // CH=5 OP=3
cfg[97] = { 1'b0, 8'h70, 8'h2}; // CH=0 OP=0
cfg[98] = { 1'b0, 8'h71, 8'h1a}; // CH=1 OP=0
cfg[99] = { 1'b0, 8'h72, 8'hfe}; // CH=2 OP=0
cfg[100] = { 1'b1, 8'h70, 8'h43}; // CH=3 OP=0
cfg[101] = { 1'b1, 8'h71, 8'hfb}; // CH=4 OP=0
cfg[102] = { 1'b1, 8'h72, 8'hfa}; // CH=5 OP=0
cfg[103] = { 1'b0, 8'h74, 8'haa}; // CH=0 OP=1
cfg[104] = { 1'b0, 8'h75, 8'h3a}; // CH=1 OP=1
cfg[105] = { 1'b0, 8'h76, 8'hfb}; // CH=2 OP=1
cfg[106] = { 1'b1, 8'h74, 8'h29}; // CH=3 OP=1
cfg[107] = { 1'b1, 8'h75, 8'hd1}; // CH=4 OP=1
cfg[108] = { 1'b1, 8'h76, 8'he6}; // CH=5 OP=1
cfg[109] = { 1'b0, 8'h78, 8'h5}; // CH=0 OP=2
cfg[110] = { 1'b0, 8'h79, 8'h3c}; // CH=1 OP=2
cfg[111] = { 1'b0, 8'h7a, 8'h7c}; // CH=2 OP=2
cfg[112] = { 1'b1, 8'h78, 8'h94}; // CH=3 OP=2
cfg[113] = { 1'b1, 8'h79, 8'h75}; // CH=4 OP=2
cfg[114] = { 1'b1, 8'h7a, 8'hd8}; // CH=5 OP=2
cfg[115] = { 1'b0, 8'h7c, 8'hbe}; // CH=0 OP=3
cfg[116] = { 1'b0, 8'h7d, 8'h61}; // CH=1 OP=3
cfg[117] = { 1'b0, 8'h7e, 8'h89}; // CH=2 OP=3
cfg[118] = { 1'b1, 8'h7c, 8'hf9}; // CH=3 OP=3
cfg[119] = { 1'b1, 8'h7d, 8'h5c}; // CH=4 OP=3
cfg[120] = { 1'b1, 8'h7e, 8'hbb}; // CH=5 OP=3
cfg[121] = { 1'b0, 8'h80, 8'ha8}; // CH=0 OP=0
cfg[122] = { 1'b0, 8'h81, 8'h99}; // CH=1 OP=0
cfg[123] = { 1'b0, 8'h82, 8'hf}; // CH=2 OP=0
cfg[124] = { 1'b1, 8'h80, 8'h95}; // CH=3 OP=0
cfg[125] = { 1'b1, 8'h81, 8'hb1}; // CH=4 OP=0
cfg[126] = { 1'b1, 8'h82, 8'heb}; // CH=5 OP=0
cfg[127] = { 1'b0, 8'h84, 8'hf1}; // CH=0 OP=1
cfg[128] = { 1'b0, 8'h85, 8'hb3}; // CH=1 OP=1
cfg[129] = { 1'b0, 8'h86, 8'h5}; // CH=2 OP=1
cfg[130] = { 1'b1, 8'h84, 8'hef}; // CH=3 OP=1
cfg[131] = { 1'b1, 8'h85, 8'hf7}; // CH=4 OP=1
cfg[132] = { 1'b1, 8'h86, 8'h0}; // CH=5 OP=1
cfg[133] = { 1'b0, 8'h88, 8'he9}; // CH=0 OP=2
cfg[134] = { 1'b0, 8'h89, 8'ha1}; // CH=1 OP=2
cfg[135] = { 1'b0, 8'h8a, 8'h3a}; // CH=2 OP=2
cfg[136] = { 1'b1, 8'h88, 8'he5}; // CH=3 OP=2
cfg[137] = { 1'b1, 8'h89, 8'hca}; // CH=4 OP=2
cfg[138] = { 1'b1, 8'h8a, 8'hb}; // CH=5 OP=2
cfg[139] = { 1'b0, 8'h8c, 8'hcb}; // CH=0 OP=3
cfg[140] = { 1'b0, 8'h8d, 8'hd0}; // CH=1 OP=3
cfg[141] = { 1'b0, 8'h8e, 8'h48}; // CH=2 OP=3
cfg[142] = { 1'b1, 8'h8c, 8'h47}; // CH=3 OP=3
cfg[143] = { 1'b1, 8'h8d, 8'h64}; // CH=4 OP=3
cfg[144] = { 1'b1, 8'h8e, 8'hbd}; // CH=5 OP=3
cfg[145] = { 1'b0, 8'h90, 8'h1f}; // CH=0 OP=0
cfg[146] = { 1'b0, 8'h91, 8'h23}; // CH=1 OP=0
cfg[147] = { 1'b0, 8'h92, 8'h1e}; // CH=2 OP=0
cfg[148] = { 1'b1, 8'h90, 8'ha8}; // CH=3 OP=0
cfg[149] = { 1'b1, 8'h91, 8'h1c}; // CH=4 OP=0
cfg[150] = { 1'b1, 8'h92, 8'h7b}; // CH=5 OP=0
cfg[151] = { 1'b0, 8'h94, 8'h64}; // CH=0 OP=1
cfg[152] = { 1'b0, 8'h95, 8'hc5}; // CH=1 OP=1
cfg[153] = { 1'b0, 8'h96, 8'h14}; // CH=2 OP=1
cfg[154] = { 1'b1, 8'h94, 8'h73}; // CH=3 OP=1
cfg[155] = { 1'b1, 8'h95, 8'h5a}; // CH=4 OP=1
cfg[156] = { 1'b1, 8'h96, 8'hc5}; // CH=5 OP=1
cfg[157] = { 1'b0, 8'h98, 8'h5e}; // CH=0 OP=2
cfg[158] = { 1'b0, 8'h99, 8'h4b}; // CH=1 OP=2
cfg[159] = { 1'b0, 8'h9a, 8'h79}; // CH=2 OP=2
cfg[160] = { 1'b1, 8'h98, 8'h63}; // CH=3 OP=2
cfg[161] = { 1'b1, 8'h99, 8'h3b}; // CH=4 OP=2
cfg[162] = { 1'b1, 8'h9a, 8'h70}; // CH=5 OP=2
cfg[163] = { 1'b0, 8'h9c, 8'h64}; // CH=0 OP=3
cfg[164] = { 1'b0, 8'h9d, 8'h24}; // CH=1 OP=3
cfg[165] = { 1'b0, 8'h9e, 8'h11}; // CH=2 OP=3
cfg[166] = { 1'b1, 8'h9c, 8'h9e}; // CH=3 OP=3
cfg[167] = { 1'b1, 8'h9d, 8'h9}; // CH=4 OP=3
cfg[168] = { 1'b1, 8'h9e, 8'hdc}; // CH=5 OP=3
cfg[169] = { 1'b0, 8'ha0, 8'haa}; // CH=0 OP=0
cfg[170] = { 1'b0, 8'ha1, 8'hd4}; // CH=1 OP=0
cfg[171] = { 1'b0, 8'ha2, 8'hac}; // CH=2 OP=0
cfg[172] = { 1'b1, 8'ha0, 8'hf2}; // CH=3 OP=0
cfg[173] = { 1'b1, 8'ha1, 8'h1b}; // CH=4 OP=0
cfg[174] = { 1'b1, 8'ha2, 8'h10}; // CH=5 OP=0
cfg[175] = { 1'b0, 8'ha4, 8'haf}; // CH=0 OP=1
cfg[176] = { 1'b0, 8'ha5, 8'h3b}; // CH=1 OP=1
cfg[177] = { 1'b0, 8'ha6, 8'h33}; // CH=2 OP=1
cfg[178] = { 1'b1, 8'ha4, 8'hcd}; // CH=3 OP=1
cfg[179] = { 1'b1, 8'ha5, 8'he3}; // CH=4 OP=1
cfg[180] = { 1'b1, 8'ha6, 8'h50}; // CH=5 OP=1
cfg[181] = { 1'b0, 8'hb0, 8'h48}; // CH=0 OP=0
cfg[182] = { 1'b0, 8'hb1, 8'h47}; // CH=1 OP=0
cfg[183] = { 1'b0, 8'hb2, 8'h15}; // CH=2 OP=0
cfg[184] = { 1'b1, 8'hb0, 8'h5c}; // CH=3 OP=0
cfg[185] = { 1'b1, 8'hb1, 8'hbb}; // CH=4 OP=0
cfg[186] = { 1'b1, 8'hb2, 8'h6f}; // CH=5 OP=0
cfg[187] = { 1'b0, 8'hb4, 8'h22}; // CH=0 OP=1
cfg[188] = { 1'b0, 8'hb5, 8'h19}; // CH=1 OP=1
cfg[189] = { 1'b0, 8'hb6, 8'hba}; // CH=2 OP=1
cfg[190] = { 1'b1, 8'hb4, 8'h9b}; // CH=3 OP=1
cfg[191] = { 1'b1, 8'hb5, 8'h7d}; // CH=4 OP=1
cfg[192] = { 1'b1, 8'hb6, 8'hf5}; // CH=5 OP=1
cfg[193] = { 1'b0, 8'hc0, 8'hb}; // CH=0 OP=0
cfg[194] = { 1'b0, 8'hc1, 8'he1}; // CH=1 OP=0
cfg[195] = { 1'b0, 8'hc2, 8'h1a}; // CH=2 OP=0
cfg[196] = { 1'b1, 8'hc0, 8'h1c}; // CH=3 OP=0
cfg[197] = { 1'b1, 8'hc1, 8'h7f}; // CH=4 OP=0
cfg[198] = { 1'b1, 8'hc2, 8'h23}; // CH=5 OP=0
cfg[199] = { 1'b0, 8'hc4, 8'hf8}; // CH=0 OP=1
cfg[200] = { 1'b0, 8'hc5, 8'h29}; // CH=1 OP=1
cfg[201] = { 1'b0, 8'hc6, 8'hf8}; // CH=2 OP=1
cfg[202] = { 1'b1, 8'hc4, 8'ha4}; // CH=3 OP=1
cfg[203] = { 1'b1, 8'hc5, 8'h1b}; // CH=4 OP=1
cfg[204] = { 1'b1, 8'hc6, 8'h13}; // CH=5 OP=1
cfg[205] = { 1'b0, 8'hd0, 8'hb5}; // CH=0 OP=0
cfg[206] = { 1'b0, 8'hd1, 8'hca}; // CH=1 OP=0
cfg[207] = { 1'b0, 8'hd2, 8'h4e}; // CH=2 OP=0
cfg[208] = { 1'b1, 8'hd0, 8'he8}; // CH=3 OP=0
cfg[209] = { 1'b1, 8'hd1, 8'h98}; // CH=4 OP=0
cfg[210] = { 1'b1, 8'hd2, 8'h32}; // CH=5 OP=0
cfg[211] = { 1'b0, 8'hd4, 8'h38}; // CH=0 OP=1
cfg[212] = { 1'b0, 8'hd5, 8'he0}; // CH=1 OP=1
cfg[213] = { 1'b0, 8'hd6, 8'h79}; // CH=2 OP=1
cfg[214] = { 1'b1, 8'hd4, 8'h4d}; // CH=3 OP=1
cfg[215] = { 1'b1, 8'hd5, 8'h3d}; // CH=4 OP=1
cfg[216] = { 1'b1, 8'hd6, 8'h34}; // CH=5 OP=1
cfg[217] = { 1'b0, 8'he0, 8'hbc}; // CH=0 OP=0
cfg[218] = { 1'b0, 8'he1, 8'h5f}; // CH=1 OP=0
cfg[219] = { 1'b0, 8'he2, 8'h4e}; // CH=2 OP=0
cfg[220] = { 1'b1, 8'he0, 8'h77}; // CH=3 OP=0
cfg[221] = { 1'b1, 8'he1, 8'hfa}; // CH=4 OP=0
cfg[222] = { 1'b1, 8'he2, 8'hcb}; // CH=5 OP=0
cfg[223] = { 1'b0, 8'he4, 8'h6c}; // CH=0 OP=1
cfg[224] = { 1'b0, 8'he5, 8'h5}; // CH=1 OP=1
cfg[225] = { 1'b0, 8'he6, 8'hac}; // CH=2 OP=1
cfg[226] = { 1'b1, 8'he4, 8'h86}; // CH=3 OP=1
cfg[227] = { 1'b1, 8'he5, 8'h21}; // CH=4 OP=1
cfg[228] = { 1'b1, 8'he6, 8'h2b}; // CH=5 OP=1
cfg[229] = { 1'b0, 8'hf0, 8'haa}; // CH=0 OP=0
cfg[230] = { 1'b0, 8'hf1, 8'h1a}; // CH=1 OP=0
cfg[231] = { 1'b0, 8'hf2, 8'h55}; // CH=2 OP=0
cfg[232] = { 1'b1, 8'hf0, 8'ha2}; // CH=3 OP=0
cfg[233] = { 1'b1, 8'hf1, 8'hbe}; // CH=4 OP=0
cfg[234] = { 1'b1, 8'hf2, 8'h70}; // CH=5 OP=0
cfg[235] = { 1'b0, 8'hf4, 8'hb5}; // CH=0 OP=1
cfg[236] = { 1'b0, 8'hf5, 8'h73}; // CH=1 OP=1
cfg[237] = { 1'b0, 8'hf6, 8'h3b}; // CH=2 OP=1
cfg[238] = { 1'b1, 8'hf4, 8'h4}; // CH=3 OP=1
cfg[239] = { 1'b1, 8'hf5, 8'h5c}; // CH=4 OP=1
cfg[240] = { 1'b1, 8'hf6, 8'hd3}; // CH=5 OP=1

cfg[241] = { 1'b0, 8'h0, 8'h00 }; // done
