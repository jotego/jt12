/* This file is part of JT12.

 
    JT12 program is free software: you can redistribute it and/or modify
    it under the terms of the GNU General Public License as published by
    the Free Software Foundation, either version 3 of the License, or
    (at your option) any later version.

    JT12 program is distributed in the hope that it will be useful,
    but WITHOUT ANY WARRANTY; without even the implied warranty of
    MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
    GNU General Public License for more details.

    You should have received a copy of the GNU General Public License
    along with JT12.  If not, see <http://www.gnu.org/licenses/>.

    Author: Jose Tejada Gomez. Twitter: @topapate
    Version: 1.0
    Date: 21-03-2019
*/

// ADPCM-A uses a LUT because it is very sensitive to rounding
// it looks like the original algorithm also used a table

module jt10_adpcma_lut(
    input              clk,        // CPU clock
    input              rst_n,
    input              cen,
    input      [8:0]   addr,       //  = {step,delta};
    output reg [11:0]  inc
);

reg [11:0] lut[0:391];

initial begin
lut[9'o00_0] = 12'o0002; lut[9'o00_1] = 12'o0006; lut[9'o00_2] = 12'o0012; lut[9'o00_3] = 12'o0016; 
lut[9'o00_4] = 12'o0022; lut[9'o00_5] = 12'o0026; lut[9'o00_6] = 12'o0032; lut[9'o00_7] = 12'o0036; 
lut[9'o01_0] = 12'o0002; lut[9'o01_1] = 12'o0006; lut[9'o01_2] = 12'o0012; lut[9'o01_3] = 12'o0016; 
lut[9'o01_4] = 12'o0023; lut[9'o01_5] = 12'o0027; lut[9'o01_6] = 12'o0033; lut[9'o01_7] = 12'o0037; 
lut[9'o02_0] = 12'o0002; lut[9'o02_1] = 12'o0007; lut[9'o02_2] = 12'o0013; lut[9'o02_3] = 12'o0020; 
lut[9'o02_4] = 12'o0025; lut[9'o02_5] = 12'o0032; lut[9'o02_6] = 12'o0036; lut[9'o02_7] = 12'o0043; 
lut[9'o03_0] = 12'o0002; lut[9'o03_1] = 12'o0007; lut[9'o03_2] = 12'o0015; lut[9'o03_3] = 12'o0022; 
lut[9'o03_4] = 12'o0027; lut[9'o03_5] = 12'o0034; lut[9'o03_6] = 12'o0042; lut[9'o03_7] = 12'o0047; 
lut[9'o04_0] = 12'o0002; lut[9'o04_1] = 12'o0010; lut[9'o04_2] = 12'o0016; lut[9'o04_3] = 12'o0024; 
lut[9'o04_4] = 12'o0031; lut[9'o04_5] = 12'o0037; lut[9'o04_6] = 12'o0045; lut[9'o04_7] = 12'o0053; 
lut[9'o05_0] = 12'o0003; lut[9'o05_1] = 12'o0011; lut[9'o05_2] = 12'o0017; lut[9'o05_3] = 12'o0025; 
lut[9'o05_4] = 12'o0034; lut[9'o05_5] = 12'o0042; lut[9'o05_6] = 12'o0050; lut[9'o05_7] = 12'o0056; 
lut[9'o06_0] = 12'o0003; lut[9'o06_1] = 12'o0012; lut[9'o06_2] = 12'o0021; lut[9'o06_3] = 12'o0030; 
lut[9'o06_4] = 12'o0037; lut[9'o06_5] = 12'o0046; lut[9'o06_6] = 12'o0055; lut[9'o06_7] = 12'o0064; 
lut[9'o07_0] = 12'o0003; lut[9'o07_1] = 12'o0013; lut[9'o07_2] = 12'o0023; lut[9'o07_3] = 12'o0033; 
lut[9'o07_4] = 12'o0042; lut[9'o07_5] = 12'o0052; lut[9'o07_6] = 12'o0062; lut[9'o07_7] = 12'o0072; 
lut[9'o10_0] = 12'o0004; lut[9'o10_1] = 12'o0014; lut[9'o10_2] = 12'o0025; lut[9'o10_3] = 12'o0035; 
lut[9'o10_4] = 12'o0046; lut[9'o10_5] = 12'o0056; lut[9'o10_6] = 12'o0067; lut[9'o10_7] = 12'o0077; 
lut[9'o11_0] = 12'o0004; lut[9'o11_1] = 12'o0015; lut[9'o11_2] = 12'o0027; lut[9'o11_3] = 12'o0040; 
lut[9'o11_4] = 12'o0051; lut[9'o11_5] = 12'o0062; lut[9'o11_6] = 12'o0074; lut[9'o11_7] = 12'o0105; 
lut[9'o12_0] = 12'o0005; lut[9'o12_1] = 12'o0017; lut[9'o12_2] = 12'o0031; lut[9'o12_3] = 12'o0043; 
lut[9'o12_4] = 12'o0056; lut[9'o12_5] = 12'o0070; lut[9'o12_6] = 12'o0102; lut[9'o12_7] = 12'o0114; 
lut[9'o13_0] = 12'o0005; lut[9'o13_1] = 12'o0020; lut[9'o13_2] = 12'o0034; lut[9'o13_3] = 12'o0047; 
lut[9'o13_4] = 12'o0062; lut[9'o13_5] = 12'o0075; lut[9'o13_6] = 12'o0111; lut[9'o13_7] = 12'o0124; 
lut[9'o14_0] = 12'o0006; lut[9'o14_1] = 12'o0022; lut[9'o14_2] = 12'o0037; lut[9'o14_3] = 12'o0053; 
lut[9'o14_4] = 12'o0070; lut[9'o14_5] = 12'o0104; lut[9'o14_6] = 12'o0121; lut[9'o14_7] = 12'o0135; 
lut[9'o15_0] = 12'o0006; lut[9'o15_1] = 12'o0024; lut[9'o15_2] = 12'o0042; lut[9'o15_3] = 12'o0060; 
lut[9'o15_4] = 12'o0075; lut[9'o15_5] = 12'o0113; lut[9'o15_6] = 12'o0131; lut[9'o15_7] = 12'o0147; 
lut[9'o16_0] = 12'o0007; lut[9'o16_1] = 12'o0026; lut[9'o16_2] = 12'o0045; lut[9'o16_3] = 12'o0064; 
lut[9'o16_4] = 12'o0103; lut[9'o16_5] = 12'o0122; lut[9'o16_6] = 12'o0141; lut[9'o16_7] = 12'o0160; 
lut[9'o17_0] = 12'o0010; lut[9'o17_1] = 12'o0030; lut[9'o17_2] = 12'o0051; lut[9'o17_3] = 12'o0071; 
lut[9'o17_4] = 12'o0112; lut[9'o17_5] = 12'o0132; lut[9'o17_6] = 12'o0153; lut[9'o17_7] = 12'o0173; 
lut[9'o20_0] = 12'o0011; lut[9'o20_1] = 12'o0033; lut[9'o20_2] = 12'o0055; lut[9'o20_3] = 12'o0077; 
lut[9'o20_4] = 12'o0122; lut[9'o20_5] = 12'o0144; lut[9'o20_6] = 12'o0166; lut[9'o20_7] = 12'o0210; 
lut[9'o21_0] = 12'o0012; lut[9'o21_1] = 12'o0036; lut[9'o21_2] = 12'o0062; lut[9'o21_3] = 12'o0106; 
lut[9'o21_4] = 12'o0132; lut[9'o21_5] = 12'o0156; lut[9'o21_6] = 12'o0202; lut[9'o21_7] = 12'o0226; 
lut[9'o22_0] = 12'o0013; lut[9'o22_1] = 12'o0041; lut[9'o22_2] = 12'o0067; lut[9'o22_3] = 12'o0115; 
lut[9'o22_4] = 12'o0143; lut[9'o22_5] = 12'o0171; lut[9'o22_6] = 12'o0217; lut[9'o22_7] = 12'o0245; 
lut[9'o23_0] = 12'o0014; lut[9'o23_1] = 12'o0044; lut[9'o23_2] = 12'o0074; lut[9'o23_3] = 12'o0124; 
lut[9'o23_4] = 12'o0155; lut[9'o23_5] = 12'o0205; lut[9'o23_6] = 12'o0235; lut[9'o23_7] = 12'o0265; 
lut[9'o24_0] = 12'o0015; lut[9'o24_1] = 12'o0050; lut[9'o24_2] = 12'o0102; lut[9'o24_3] = 12'o0135; 
lut[9'o24_4] = 12'o0170; lut[9'o24_5] = 12'o0223; lut[9'o24_6] = 12'o0255; lut[9'o24_7] = 12'o0310; 
lut[9'o25_0] = 12'o0016; lut[9'o25_1] = 12'o0054; lut[9'o25_2] = 12'o0111; lut[9'o25_3] = 12'o0147; 
lut[9'o25_4] = 12'o0204; lut[9'o25_5] = 12'o0242; lut[9'o25_6] = 12'o0277; lut[9'o25_7] = 12'o0335; 
lut[9'o26_0] = 12'o0020; lut[9'o26_1] = 12'o0060; lut[9'o26_2] = 12'o0121; lut[9'o26_3] = 12'o0161; 
lut[9'o26_4] = 12'o0222; lut[9'o26_5] = 12'o0262; lut[9'o26_6] = 12'o0323; lut[9'o26_7] = 12'o0363; 
lut[9'o27_0] = 12'o0021; lut[9'o27_1] = 12'o0065; lut[9'o27_2] = 12'o0131; lut[9'o27_3] = 12'o0175; 
lut[9'o27_4] = 12'o0240; lut[9'o27_5] = 12'o0304; lut[9'o27_6] = 12'o0350; lut[9'o27_7] = 12'o0414; 
lut[9'o30_0] = 12'o0023; lut[9'o30_1] = 12'o0072; lut[9'o30_2] = 12'o0142; lut[9'o30_3] = 12'o0211; 
lut[9'o30_4] = 12'o0260; lut[9'o30_5] = 12'o0327; lut[9'o30_6] = 12'o0377; lut[9'o30_7] = 12'o0446; 
lut[9'o31_0] = 12'o0025; lut[9'o31_1] = 12'o0100; lut[9'o31_2] = 12'o0154; lut[9'o31_3] = 12'o0227; 
lut[9'o31_4] = 12'o0302; lut[9'o31_5] = 12'o0355; lut[9'o31_6] = 12'o0431; lut[9'o31_7] = 12'o0504; 
lut[9'o32_0] = 12'o0027; lut[9'o32_1] = 12'o0107; lut[9'o32_2] = 12'o0166; lut[9'o32_3] = 12'o0246; 
lut[9'o32_4] = 12'o0325; lut[9'o32_5] = 12'o0405; lut[9'o32_6] = 12'o0464; lut[9'o32_7] = 12'o0544; 
lut[9'o33_0] = 12'o0032; lut[9'o33_1] = 12'o0116; lut[9'o33_2] = 12'o0202; lut[9'o33_3] = 12'o0266; 
lut[9'o33_4] = 12'o0353; lut[9'o33_5] = 12'o0437; lut[9'o33_6] = 12'o0523; lut[9'o33_7] = 12'o0607; 
lut[9'o34_0] = 12'o0034; lut[9'o34_1] = 12'o0126; lut[9'o34_2] = 12'o0217; lut[9'o34_3] = 12'o0311; 
lut[9'o34_4] = 12'o0402; lut[9'o34_5] = 12'o0474; lut[9'o34_6] = 12'o0565; lut[9'o34_7] = 12'o0657; 
lut[9'o35_0] = 12'o0037; lut[9'o35_1] = 12'o0136; lut[9'o35_2] = 12'o0236; lut[9'o35_3] = 12'o0335; 
lut[9'o35_4] = 12'o0434; lut[9'o35_5] = 12'o0533; lut[9'o35_6] = 12'o0633; lut[9'o35_7] = 12'o0732; 
lut[9'o36_0] = 12'o0042; lut[9'o36_1] = 12'o0150; lut[9'o36_2] = 12'o0256; lut[9'o36_3] = 12'o0364; 
lut[9'o36_4] = 12'o0471; lut[9'o36_5] = 12'o0577; lut[9'o36_6] = 12'o0705; lut[9'o36_7] = 12'o1013; 
lut[9'o37_0] = 12'o0046; lut[9'o37_1] = 12'o0163; lut[9'o37_2] = 12'o0277; lut[9'o37_3] = 12'o0414; 
lut[9'o37_4] = 12'o0531; lut[9'o37_5] = 12'o0646; lut[9'o37_6] = 12'o0762; lut[9'o37_7] = 12'o1077; 
lut[9'o40_0] = 12'o0052; lut[9'o40_1] = 12'o0176; lut[9'o40_2] = 12'o0322; lut[9'o40_3] = 12'o0446; 
lut[9'o40_4] = 12'o0573; lut[9'o40_5] = 12'o0717; lut[9'o40_6] = 12'o1043; lut[9'o40_7] = 12'o1167; 
lut[9'o41_0] = 12'o0056; lut[9'o41_1] = 12'o0213; lut[9'o41_2] = 12'o0347; lut[9'o41_3] = 12'o0504; 
lut[9'o41_4] = 12'o0641; lut[9'o41_5] = 12'o0776; lut[9'o41_6] = 12'o1132; lut[9'o41_7] = 12'o1267; 
lut[9'o42_0] = 12'o0063; lut[9'o42_1] = 12'o0231; lut[9'o42_2] = 12'o0377; lut[9'o42_3] = 12'o0545; 
lut[9'o42_4] = 12'o0713; lut[9'o42_5] = 12'o1061; lut[9'o42_6] = 12'o1227; lut[9'o42_7] = 12'o1375; 
lut[9'o43_0] = 12'o0070; lut[9'o43_1] = 12'o0250; lut[9'o43_2] = 12'o0430; lut[9'o43_3] = 12'o0610; 
lut[9'o43_4] = 12'o0771; lut[9'o43_5] = 12'o1151; lut[9'o43_6] = 12'o1331; lut[9'o43_7] = 12'o1511; 
lut[9'o44_0] = 12'o0075; lut[9'o44_1] = 12'o0271; lut[9'o44_2] = 12'o0464; lut[9'o44_3] = 12'o0660; 
lut[9'o44_4] = 12'o1053; lut[9'o44_5] = 12'o1247; lut[9'o44_6] = 12'o1442; lut[9'o44_7] = 12'o1636; 
lut[9'o45_0] = 12'o0104; lut[9'o45_1] = 12'o0314; lut[9'o45_2] = 12'o0524; lut[9'o45_3] = 12'o0734; 
lut[9'o45_4] = 12'o1144; lut[9'o45_5] = 12'o1354; lut[9'o45_6] = 12'o1564; lut[9'o45_7] = 12'o1774; 
lut[9'o46_0] = 12'o0112; lut[9'o46_1] = 12'o0340; lut[9'o46_2] = 12'o0565; lut[9'o46_3] = 12'o1013; 
lut[9'o46_4] = 12'o1240; lut[9'o46_5] = 12'o1466; lut[9'o46_6] = 12'o1713; lut[9'o46_7] = 12'o2141; 
lut[9'o47_0] = 12'o0122; lut[9'o47_1] = 12'o0366; lut[9'o47_2] = 12'o0633; lut[9'o47_3] = 12'o1077; 
lut[9'o47_4] = 12'o1344; lut[9'o47_5] = 12'o1610; lut[9'o47_6] = 12'o2055; lut[9'o47_7] = 12'o2321; 
lut[9'o50_0] = 12'o0132; lut[9'o50_1] = 12'o0417; lut[9'o50_2] = 12'o0704; lut[9'o50_3] = 12'o1171; 
lut[9'o50_4] = 12'o1456; lut[9'o50_5] = 12'o1743; lut[9'o50_6] = 12'o2230; lut[9'o50_7] = 12'o2515; 
lut[9'o51_0] = 12'o0143; lut[9'o51_1] = 12'o0452; lut[9'o51_2] = 12'o0761; lut[9'o51_3] = 12'o1270; 
lut[9'o51_4] = 12'o1577; lut[9'o51_5] = 12'o2106; lut[9'o51_6] = 12'o2415; lut[9'o51_7] = 12'o2724; 
lut[9'o52_0] = 12'o0155; lut[9'o52_1] = 12'o0510; lut[9'o52_2] = 12'o1043; lut[9'o52_3] = 12'o1376; 
lut[9'o52_4] = 12'o1731; lut[9'o52_5] = 12'o2264; lut[9'o52_6] = 12'o2617; lut[9'o52_7] = 12'o3152; 
lut[9'o53_0] = 12'o0170; lut[9'o53_1] = 12'o0551; lut[9'o53_2] = 12'o1131; lut[9'o53_3] = 12'o1512; 
lut[9'o53_4] = 12'o2073; lut[9'o53_5] = 12'o2454; lut[9'o53_6] = 12'o3034; lut[9'o53_7] = 12'o3415; 
lut[9'o54_0] = 12'o0204; lut[9'o54_1] = 12'o0615; lut[9'o54_2] = 12'o1226; lut[9'o54_3] = 12'o1637; 
lut[9'o54_4] = 12'o2250; lut[9'o54_5] = 12'o2661; lut[9'o54_6] = 12'o3272; lut[9'o54_7] = 12'o3703; 
lut[9'o55_0] = 12'o0221; lut[9'o55_1] = 12'o0665; lut[9'o55_2] = 12'o1330; lut[9'o55_3] = 12'o1774;// Not sure if these should clip at 11 bits or not
lut[9'o55_4] = 12'o2437; lut[9'o55_5] = 12'o3103; lut[9'o55_6] = 12'o3546; lut[9'o55_7] = 12'o4212;//12'o3777; 
lut[9'o56_0] = 12'o0240; lut[9'o56_1] = 12'o0740; lut[9'o56_2] = 12'o1441; lut[9'o56_3] = 12'o2141; 
lut[9'o56_4] = 12'o2642; lut[9'o56_5] = 12'o3342; lut[9'o56_6] = 12'o4043; lut[9'o56_7] = 12'o4543;//12'o3777; lut[9'o56_7] = 12'o3777; 
lut[9'o57_0] = 12'o0260; lut[9'o57_1] = 12'o1021; lut[9'o57_2] = 12'o1561; lut[9'o57_3] = 12'o2322; 
lut[9'o57_4] = 12'o3063; lut[9'o57_5] = 12'o3624; lut[9'o57_6] = 12'o4364; lut[9'o57_7] = 12'o5125;//12'o3777; lut[9'o57_7] = 12'o3777;  
lut[9'o60_0] = 12'o0302; lut[9'o60_1] = 12'o1106; lut[9'o60_2] = 12'o1712; lut[9'o60_3] = 12'o2516; 
lut[9'o60_4] = 12'o3322; lut[9'o60_5] = 12'o4126; lut[9'o60_6] = 12'o4732; lut[9'o60_7] = 12'o5536;//12'o3777; lut[9'o60_6] = 12'o3777; lut[9'o60_7] = 12'o3777; 
end

always @(posedge clk or negedge rst_n) 
    if(!rst_n)
        inc <= 'd0;
    else if(cen)
        inc <= lut[addr];

endmodule // jt10_adpcma_lut
