cfg[0] = { 1'b0, 8'ha0, 8'h0};
cfg[1] = { 1'b0, 8'ha4, 8'h24};
cfg[2] = { 1'b0, 8'hb0, 8'h7};
cfg[3] = { 1'b0, 8'hb4, 8'h0};
cfg[4] = { 1'b0, 8'h30, 8'h1};
cfg[5] = { 1'b0, 8'h40, 8'h7f};
cfg[6] = { 1'b0, 8'h50, 8'h1f};
cfg[7] = { 1'b0, 8'h60, 8'h14};
cfg[8] = { 1'b0, 8'h70, 8'he};
cfg[9] = { 1'b0, 8'h80, 8'haf};
cfg[10] = { 1'b0, 8'h90, 8'h0};
cfg[11] = { 1'b0, 8'h38, 8'h1};
cfg[12] = { 1'b0, 8'h48, 8'h7f};
cfg[13] = { 1'b0, 8'h58, 8'h1f};
cfg[14] = { 1'b0, 8'h68, 8'h14};
cfg[15] = { 1'b0, 8'h78, 8'he};
cfg[16] = { 1'b0, 8'h88, 8'haf};
cfg[17] = { 1'b0, 8'h98, 8'h0};
cfg[18] = { 1'b0, 8'h34, 8'h1};
cfg[19] = { 1'b0, 8'h44, 8'h7f};
cfg[20] = { 1'b0, 8'h54, 8'h1f};
cfg[21] = { 1'b0, 8'h64, 8'h14};
cfg[22] = { 1'b0, 8'h74, 8'he};
cfg[23] = { 1'b0, 8'h84, 8'haf};
cfg[24] = { 1'b0, 8'h94, 8'h0};
cfg[25] = { 1'b0, 8'h3c, 8'h1};
cfg[26] = { 1'b0, 8'h4c, 8'h7f};
cfg[27] = { 1'b0, 8'h5c, 8'h1f};
cfg[28] = { 1'b0, 8'h6c, 8'h14};
cfg[29] = { 1'b0, 8'h7c, 8'he};
cfg[30] = { 1'b0, 8'h8c, 8'haf};
cfg[31] = { 1'b0, 8'h9c, 8'h0};
cfg[32] = { 1'b0, 8'ha1, 8'h0};
cfg[33] = { 1'b0, 8'ha5, 8'h24};
cfg[34] = { 1'b0, 8'hb1, 8'h7};
cfg[35] = { 1'b0, 8'hb5, 8'h0};
cfg[36] = { 1'b0, 8'h31, 8'h1};
cfg[37] = { 1'b0, 8'h41, 8'h7f};
cfg[38] = { 1'b0, 8'h51, 8'h1f};
cfg[39] = { 1'b0, 8'h61, 8'h14};
cfg[40] = { 1'b0, 8'h71, 8'he};
cfg[41] = { 1'b0, 8'h81, 8'haf};
cfg[42] = { 1'b0, 8'h91, 8'h0};
cfg[43] = { 1'b0, 8'h39, 8'h1};
cfg[44] = { 1'b0, 8'h49, 8'h7f};
cfg[45] = { 1'b0, 8'h59, 8'h1f};
cfg[46] = { 1'b0, 8'h69, 8'h14};
cfg[47] = { 1'b0, 8'h79, 8'he};
cfg[48] = { 1'b0, 8'h89, 8'haf};
cfg[49] = { 1'b0, 8'h99, 8'h0};
cfg[50] = { 1'b0, 8'h35, 8'h1};
cfg[51] = { 1'b0, 8'h45, 8'h7f};
cfg[52] = { 1'b0, 8'h55, 8'h1f};
cfg[53] = { 1'b0, 8'h65, 8'h14};
cfg[54] = { 1'b0, 8'h75, 8'he};
cfg[55] = { 1'b0, 8'h85, 8'haf};
cfg[56] = { 1'b0, 8'h95, 8'h0};
cfg[57] = { 1'b0, 8'h3d, 8'h1};
cfg[58] = { 1'b0, 8'h4d, 8'h7f};
cfg[59] = { 1'b0, 8'h5d, 8'h1f};
cfg[60] = { 1'b0, 8'h6d, 8'h14};
cfg[61] = { 1'b0, 8'h7d, 8'he};
cfg[62] = { 1'b0, 8'h8d, 8'haf};
cfg[63] = { 1'b0, 8'h9d, 8'h0};
cfg[64] = { 1'b0, 8'ha2, 8'h0};
cfg[65] = { 1'b0, 8'ha6, 8'h24};
cfg[66] = { 1'b0, 8'hb2, 8'h7};
cfg[67] = { 1'b0, 8'hb6, 8'h0};
cfg[68] = { 1'b0, 8'h32, 8'h1};
cfg[69] = { 1'b0, 8'h42, 8'h7f};
cfg[70] = { 1'b0, 8'h52, 8'h1f};
cfg[71] = { 1'b0, 8'h62, 8'h14};
cfg[72] = { 1'b0, 8'h72, 8'he};
cfg[73] = { 1'b0, 8'h82, 8'haf};
cfg[74] = { 1'b0, 8'h92, 8'h0};
cfg[75] = { 1'b0, 8'h3a, 8'h1};
cfg[76] = { 1'b0, 8'h4a, 8'h7f};
cfg[77] = { 1'b0, 8'h5a, 8'h1f};
cfg[78] = { 1'b0, 8'h6a, 8'h14};
cfg[79] = { 1'b0, 8'h7a, 8'he};
cfg[80] = { 1'b0, 8'h8a, 8'haf};
cfg[81] = { 1'b0, 8'h9a, 8'h0};
cfg[82] = { 1'b0, 8'h36, 8'h1};
cfg[83] = { 1'b0, 8'h46, 8'h7f};
cfg[84] = { 1'b0, 8'h56, 8'h1f};
cfg[85] = { 1'b0, 8'h66, 8'h14};
cfg[86] = { 1'b0, 8'h76, 8'he};
cfg[87] = { 1'b0, 8'h86, 8'haf};
cfg[88] = { 1'b0, 8'h96, 8'h0};
cfg[89] = { 1'b0, 8'h3e, 8'h1};
cfg[90] = { 1'b0, 8'h4e, 8'h7f};
cfg[91] = { 1'b0, 8'h5e, 8'h1f};
cfg[92] = { 1'b0, 8'h6e, 8'h14};
cfg[93] = { 1'b0, 8'h7e, 8'he};
cfg[94] = { 1'b0, 8'h8e, 8'haf};
cfg[95] = { 1'b0, 8'h9e, 8'h0};
cfg[96] = { 1'b1, 8'ha0, 8'h0};
cfg[97] = { 1'b1, 8'ha4, 8'h24};
cfg[98] = { 1'b1, 8'hb0, 8'h7};
cfg[99] = { 1'b1, 8'hb4, 8'h0};
cfg[100] = { 1'b1, 8'h30, 8'h1};
cfg[101] = { 1'b1, 8'h40, 8'h7f};
cfg[102] = { 1'b1, 8'h50, 8'h1f};
cfg[103] = { 1'b1, 8'h60, 8'h14};
cfg[104] = { 1'b1, 8'h70, 8'he};
cfg[105] = { 1'b1, 8'h80, 8'haf};
cfg[106] = { 1'b1, 8'h90, 8'h0};
cfg[107] = { 1'b1, 8'h38, 8'h1};
cfg[108] = { 1'b1, 8'h48, 8'h7f};
cfg[109] = { 1'b1, 8'h58, 8'h1f};
cfg[110] = { 1'b1, 8'h68, 8'h14};
cfg[111] = { 1'b1, 8'h78, 8'he};
cfg[112] = { 1'b1, 8'h88, 8'haf};
cfg[113] = { 1'b1, 8'h98, 8'h0};
cfg[114] = { 1'b1, 8'h34, 8'h1};
cfg[115] = { 1'b1, 8'h44, 8'h7f};
cfg[116] = { 1'b1, 8'h54, 8'h1f};
cfg[117] = { 1'b1, 8'h64, 8'h14};
cfg[118] = { 1'b1, 8'h74, 8'he};
cfg[119] = { 1'b1, 8'h84, 8'haf};
cfg[120] = { 1'b1, 8'h94, 8'h0};
cfg[121] = { 1'b1, 8'h3c, 8'h1};
cfg[122] = { 1'b1, 8'h4c, 8'h7f};
cfg[123] = { 1'b1, 8'h5c, 8'h1f};
cfg[124] = { 1'b1, 8'h6c, 8'h14};
cfg[125] = { 1'b1, 8'h7c, 8'he};
cfg[126] = { 1'b1, 8'h8c, 8'haf};
cfg[127] = { 1'b1, 8'h9c, 8'h0};
cfg[128] = { 1'b1, 8'ha1, 8'h0};
cfg[129] = { 1'b1, 8'ha5, 8'h24};
cfg[130] = { 1'b1, 8'hb1, 8'h7};
cfg[131] = { 1'b1, 8'hb5, 8'h0};
cfg[132] = { 1'b1, 8'h31, 8'h1};
cfg[133] = { 1'b1, 8'h41, 8'h7f};
cfg[134] = { 1'b1, 8'h51, 8'h1f};
cfg[135] = { 1'b1, 8'h61, 8'h14};
cfg[136] = { 1'b1, 8'h71, 8'he};
cfg[137] = { 1'b1, 8'h81, 8'haf};
cfg[138] = { 1'b1, 8'h91, 8'h0};
cfg[139] = { 1'b1, 8'h39, 8'h1};
cfg[140] = { 1'b1, 8'h49, 8'h7f};
cfg[141] = { 1'b1, 8'h59, 8'h1f};
cfg[142] = { 1'b1, 8'h69, 8'h14};
cfg[143] = { 1'b1, 8'h79, 8'he};
cfg[144] = { 1'b1, 8'h89, 8'haf};
cfg[145] = { 1'b1, 8'h99, 8'h0};
cfg[146] = { 1'b1, 8'h35, 8'h1};
cfg[147] = { 1'b1, 8'h45, 8'h7f};
cfg[148] = { 1'b1, 8'h55, 8'h1f};
cfg[149] = { 1'b1, 8'h65, 8'h14};
cfg[150] = { 1'b1, 8'h75, 8'he};
cfg[151] = { 1'b1, 8'h85, 8'haf};
cfg[152] = { 1'b1, 8'h95, 8'h0};
cfg[153] = { 1'b1, 8'h3d, 8'h1};
cfg[154] = { 1'b1, 8'h4d, 8'h7f};
cfg[155] = { 1'b1, 8'h5d, 8'h1f};
cfg[156] = { 1'b1, 8'h6d, 8'h14};
cfg[157] = { 1'b1, 8'h7d, 8'he};
cfg[158] = { 1'b1, 8'h8d, 8'haf};
cfg[159] = { 1'b1, 8'h9d, 8'h0};
cfg[160] = { 1'b1, 8'ha2, 8'h0};
cfg[161] = { 1'b1, 8'ha6, 8'h24};
cfg[162] = { 1'b1, 8'hb2, 8'h7};
cfg[163] = { 1'b1, 8'hb6, 8'h0};
cfg[164] = { 1'b1, 8'h32, 8'h1};
cfg[165] = { 1'b1, 8'h42, 8'h7f};
cfg[166] = { 1'b1, 8'h52, 8'h1f};
cfg[167] = { 1'b1, 8'h62, 8'h14};
cfg[168] = { 1'b1, 8'h72, 8'he};
cfg[169] = { 1'b1, 8'h82, 8'haf};
cfg[170] = { 1'b1, 8'h92, 8'h0};
cfg[171] = { 1'b1, 8'h3a, 8'h1};
cfg[172] = { 1'b1, 8'h4a, 8'h7f};
cfg[173] = { 1'b1, 8'h5a, 8'h1f};
cfg[174] = { 1'b1, 8'h6a, 8'h14};
cfg[175] = { 1'b1, 8'h7a, 8'he};
cfg[176] = { 1'b1, 8'h8a, 8'haf};
cfg[177] = { 1'b1, 8'h9a, 8'h0};
cfg[178] = { 1'b1, 8'h36, 8'h1};
cfg[179] = { 1'b1, 8'h46, 8'h7f};
cfg[180] = { 1'b1, 8'h56, 8'h1f};
cfg[181] = { 1'b1, 8'h66, 8'h14};
cfg[182] = { 1'b1, 8'h76, 8'he};
cfg[183] = { 1'b1, 8'h86, 8'haf};
cfg[184] = { 1'b1, 8'h96, 8'h0};
cfg[185] = { 1'b1, 8'h3e, 8'h1};
cfg[186] = { 1'b1, 8'h4e, 8'h7f};
cfg[187] = { 1'b1, 8'h5e, 8'h1f};
cfg[188] = { 1'b1, 8'h6e, 8'h14};
cfg[189] = { 1'b1, 8'h7e, 8'he};
cfg[190] = { 1'b1, 8'h8e, 8'haf};
cfg[191] = { 1'b1, 8'h9e, 8'h0};
cfg[192] = { 1'b0, 8'h28, 8'hf0};
cfg[193] = { 1'b0, 8'h28, 8'hf1};
cfg[194] = { 1'b0, 8'h28, 8'hf2};
cfg[195] = { 1'b0, 8'h28, 8'hf4};
cfg[196] = { 1'b0, 8'h28, 8'hf5};
cfg[197] = { 1'b0, 8'h28, 8'hf6};
cfg[198] = { 1'b0, 8'h1, 8'hff};
cfg[199] = { 1'b0, 8'h28, 8'h0};
cfg[200] = { 1'b0, 8'h28, 8'h1};
cfg[201] = { 1'b0, 8'h28, 8'h2};
cfg[202] = { 1'b0, 8'h28, 8'h4};
cfg[203] = { 1'b0, 8'h28, 8'h5};
cfg[204] = { 1'b0, 8'h28, 8'h6};
cfg[205] = { 1'b0, 8'h1, 8'hff};
cfg[206] = { 1'b0, 8'h40, 8'h0};
cfg[207] = { 1'b0, 8'h50, 8'h12};
cfg[208] = { 1'b0, 8'ha4, 8'hf};
cfg[209] = { 1'b0, 8'hb0, 8'h7};
cfg[210] = { 1'b0, 8'hb4, 8'hc0};
cfg[211] = { 1'b0, 8'h60, 8'h12};
cfg[212] = { 1'b0, 8'h70, 8'h12};
cfg[213] = { 1'b0, 8'h80, 8'h4f};
cfg[214] = { 1'b0, 8'h28, 8'h10};
cfg[215] = { 1'b0, 8'h1, 8'hff};
cfg[216] = { 1'b0, 8'h1, 8'hff};
cfg[217] = { 1'b0, 8'h1, 8'hff};
cfg[218] = { 1'b0, 8'h28, 8'h10};
cfg[219] = { 1'b0, 8'h1, 8'hff};
cfg[220] = { 1'b0, 8'h1, 8'hff};
cfg[221] = { 1'b0, 8'h1, 8'hff};
cfg[222] = { 1'b0, 8'h28, 8'h0};
cfg[223] = { 1'b0, 8'h1, 8'hff};
cfg[224] = { 1'b0, 8'h1, 8'hff};
cfg[225] = { 1'b0, 8'h1, 8'hff};
cfg[226] = { 1'b0, 8'h28, 8'h10};
cfg[227] = { 1'b0, 8'h1, 8'hff};
cfg[228] = { 1'b0, 8'h1, 8'hff};
cfg[229] = { 1'b0, 8'h1, 8'hff};
cfg[230] = { 1'b0, 8'h28, 8'h0};
cfg[231] = { 1'b0, 8'h1, 8'hff};
cfg[232] = { 1'b0, 8'h1, 8'hff};
cfg[233] = { 1'b0, 8'h1, 8'hff};
cfg[234] = { 1'b0, 8'h50, 8'h1f};
cfg[235] = { 1'b0, 8'h28, 8'h10};
cfg[236] = { 1'b0, 8'h1, 8'hff};
cfg[237] = { 1'b0, 8'h1, 8'hff};
cfg[238] = { 1'b0, 8'h1, 8'hff};
cfg[239] = { 1'b0, 8'h28, 8'h10};
cfg[240] = { 1'b0, 8'h1, 8'hff};
cfg[241] = { 1'b0, 8'h1, 8'hff};
cfg[242] = { 1'b0, 8'h1, 8'hff};
cfg[243] = { 1'b0, 8'h28, 8'h0};
cfg[244] = { 1'b0, 8'h1, 8'hff};
cfg[245] = { 1'b0, 8'h60, 8'h0};
cfg[246] = { 1'b0, 8'h70, 8'h0};
cfg[247] = { 1'b0, 8'h80, 8'h0};
cfg[248] = { 1'b0, 8'h28, 8'h10};
cfg[249] = { 1'b0, 8'h1, 8'hff};
cfg[250] = { 1'b0, 8'h28, 8'h0};
cfg[251] = { 1'b0, 8'h1, 8'hff};
cfg[252] = { 1'b0, 8'h28, 8'h10};
cfg[253] = { 1'b0, 8'h1, 8'hff};
cfg[254] = { 1'b0, 8'h1, 8'hff};
cfg[255] = { 1'b0, 8'h1, 8'hff};
cfg[256] = { 1'b0, 8'h28, 8'h0};
cfg[257] = { 1'b0, 8'h1, 8'hff};

cfg[258] = { 1'b0, 8'h0, 8'h00 }; // done
