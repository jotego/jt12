cfg[0] = { 1'b0, 8'ha0, 8'h0};
cfg[1] = { 1'b0, 8'ha4, 8'h24};
cfg[2] = { 1'b0, 8'hb0, 8'h7};
cfg[3] = { 1'b0, 8'hb4, 8'h0};
cfg[4] = { 1'b0, 8'h30, 8'h1};
cfg[5] = { 1'b0, 8'h40, 8'h7f};
cfg[6] = { 1'b0, 8'h50, 8'h1f};
cfg[7] = { 1'b0, 8'h60, 8'h14};
cfg[8] = { 1'b0, 8'h70, 8'he};
cfg[9] = { 1'b0, 8'h80, 8'haf};
cfg[10] = { 1'b0, 8'h90, 8'h0};
cfg[11] = { 1'b0, 8'h38, 8'h1};
cfg[12] = { 1'b0, 8'h48, 8'h7f};
cfg[13] = { 1'b0, 8'h58, 8'h1f};
cfg[14] = { 1'b0, 8'h68, 8'h14};
cfg[15] = { 1'b0, 8'h78, 8'he};
cfg[16] = { 1'b0, 8'h88, 8'haf};
cfg[17] = { 1'b0, 8'h98, 8'h0};
cfg[18] = { 1'b0, 8'h34, 8'h1};
cfg[19] = { 1'b0, 8'h44, 8'h7f};
cfg[20] = { 1'b0, 8'h54, 8'h1f};
cfg[21] = { 1'b0, 8'h64, 8'h14};
cfg[22] = { 1'b0, 8'h74, 8'he};
cfg[23] = { 1'b0, 8'h84, 8'haf};
cfg[24] = { 1'b0, 8'h94, 8'h0};
cfg[25] = { 1'b0, 8'h3c, 8'h1};
cfg[26] = { 1'b0, 8'h4c, 8'h7f};
cfg[27] = { 1'b0, 8'h5c, 8'h1f};
cfg[28] = { 1'b0, 8'h6c, 8'h14};
cfg[29] = { 1'b0, 8'h7c, 8'he};
cfg[30] = { 1'b0, 8'h8c, 8'haf};
cfg[31] = { 1'b0, 8'h9c, 8'h0};
cfg[32] = { 1'b0, 8'ha1, 8'h0};
cfg[33] = { 1'b0, 8'ha5, 8'h24};
cfg[34] = { 1'b0, 8'hb1, 8'h7};
cfg[35] = { 1'b0, 8'hb5, 8'h0};
cfg[36] = { 1'b0, 8'h31, 8'h1};
cfg[37] = { 1'b0, 8'h41, 8'h7f};
cfg[38] = { 1'b0, 8'h51, 8'h1f};
cfg[39] = { 1'b0, 8'h61, 8'h14};
cfg[40] = { 1'b0, 8'h71, 8'he};
cfg[41] = { 1'b0, 8'h81, 8'haf};
cfg[42] = { 1'b0, 8'h91, 8'h0};
cfg[43] = { 1'b0, 8'h39, 8'h1};
cfg[44] = { 1'b0, 8'h49, 8'h7f};
cfg[45] = { 1'b0, 8'h59, 8'h1f};
cfg[46] = { 1'b0, 8'h69, 8'h14};
cfg[47] = { 1'b0, 8'h79, 8'he};
cfg[48] = { 1'b0, 8'h89, 8'haf};
cfg[49] = { 1'b0, 8'h99, 8'h0};
cfg[50] = { 1'b0, 8'h35, 8'h1};
cfg[51] = { 1'b0, 8'h45, 8'h7f};
cfg[52] = { 1'b0, 8'h55, 8'h1f};
cfg[53] = { 1'b0, 8'h65, 8'h14};
cfg[54] = { 1'b0, 8'h75, 8'he};
cfg[55] = { 1'b0, 8'h85, 8'haf};
cfg[56] = { 1'b0, 8'h95, 8'h0};
cfg[57] = { 1'b0, 8'h3d, 8'h1};
cfg[58] = { 1'b0, 8'h4d, 8'h7f};
cfg[59] = { 1'b0, 8'h5d, 8'h1f};
cfg[60] = { 1'b0, 8'h6d, 8'h14};
cfg[61] = { 1'b0, 8'h7d, 8'he};
cfg[62] = { 1'b0, 8'h8d, 8'haf};
cfg[63] = { 1'b0, 8'h9d, 8'h0};
cfg[64] = { 1'b0, 8'ha2, 8'h0};
cfg[65] = { 1'b0, 8'ha6, 8'h24};
cfg[66] = { 1'b0, 8'hb2, 8'h7};
cfg[67] = { 1'b0, 8'hb6, 8'h0};
cfg[68] = { 1'b0, 8'h32, 8'h1};
cfg[69] = { 1'b0, 8'h42, 8'h7f};
cfg[70] = { 1'b0, 8'h52, 8'h1f};
cfg[71] = { 1'b0, 8'h62, 8'h14};
cfg[72] = { 1'b0, 8'h72, 8'he};
cfg[73] = { 1'b0, 8'h82, 8'haf};
cfg[74] = { 1'b0, 8'h92, 8'h0};
cfg[75] = { 1'b0, 8'h3a, 8'h1};
cfg[76] = { 1'b0, 8'h4a, 8'h7f};
cfg[77] = { 1'b0, 8'h5a, 8'h1f};
cfg[78] = { 1'b0, 8'h6a, 8'h14};
cfg[79] = { 1'b0, 8'h7a, 8'he};
cfg[80] = { 1'b0, 8'h8a, 8'haf};
cfg[81] = { 1'b0, 8'h9a, 8'h0};
cfg[82] = { 1'b0, 8'h36, 8'h1};
cfg[83] = { 1'b0, 8'h46, 8'h7f};
cfg[84] = { 1'b0, 8'h56, 8'h1f};
cfg[85] = { 1'b0, 8'h66, 8'h14};
cfg[86] = { 1'b0, 8'h76, 8'he};
cfg[87] = { 1'b0, 8'h86, 8'haf};
cfg[88] = { 1'b0, 8'h96, 8'h0};
cfg[89] = { 1'b0, 8'h3e, 8'h1};
cfg[90] = { 1'b0, 8'h4e, 8'h7f};
cfg[91] = { 1'b0, 8'h5e, 8'h1f};
cfg[92] = { 1'b0, 8'h6e, 8'h14};
cfg[93] = { 1'b0, 8'h7e, 8'he};
cfg[94] = { 1'b0, 8'h8e, 8'haf};
cfg[95] = { 1'b0, 8'h9e, 8'h0};
cfg[96] = { 1'b1, 8'ha0, 8'h0};
cfg[97] = { 1'b1, 8'ha4, 8'h24};
cfg[98] = { 1'b1, 8'hb0, 8'h7};
cfg[99] = { 1'b1, 8'hb4, 8'h0};
cfg[100] = { 1'b1, 8'h30, 8'h1};
cfg[101] = { 1'b1, 8'h40, 8'h7f};
cfg[102] = { 1'b1, 8'h50, 8'h1f};
cfg[103] = { 1'b1, 8'h60, 8'h14};
cfg[104] = { 1'b1, 8'h70, 8'he};
cfg[105] = { 1'b1, 8'h80, 8'haf};
cfg[106] = { 1'b1, 8'h90, 8'h0};
cfg[107] = { 1'b1, 8'h38, 8'h1};
cfg[108] = { 1'b1, 8'h48, 8'h7f};
cfg[109] = { 1'b1, 8'h58, 8'h1f};
cfg[110] = { 1'b1, 8'h68, 8'h14};
cfg[111] = { 1'b1, 8'h78, 8'he};
cfg[112] = { 1'b1, 8'h88, 8'haf};
cfg[113] = { 1'b1, 8'h98, 8'h0};
cfg[114] = { 1'b1, 8'h34, 8'h1};
cfg[115] = { 1'b1, 8'h44, 8'h7f};
cfg[116] = { 1'b1, 8'h54, 8'h1f};
cfg[117] = { 1'b1, 8'h64, 8'h14};
cfg[118] = { 1'b1, 8'h74, 8'he};
cfg[119] = { 1'b1, 8'h84, 8'haf};
cfg[120] = { 1'b1, 8'h94, 8'h0};
cfg[121] = { 1'b1, 8'h3c, 8'h1};
cfg[122] = { 1'b1, 8'h4c, 8'h7f};
cfg[123] = { 1'b1, 8'h5c, 8'h1f};
cfg[124] = { 1'b1, 8'h6c, 8'h14};
cfg[125] = { 1'b1, 8'h7c, 8'he};
cfg[126] = { 1'b1, 8'h8c, 8'haf};
cfg[127] = { 1'b1, 8'h9c, 8'h0};
cfg[128] = { 1'b1, 8'ha1, 8'h0};
cfg[129] = { 1'b1, 8'ha5, 8'h24};
cfg[130] = { 1'b1, 8'hb1, 8'h7};
cfg[131] = { 1'b1, 8'hb5, 8'h0};
cfg[132] = { 1'b1, 8'h31, 8'h1};
cfg[133] = { 1'b1, 8'h41, 8'h7f};
cfg[134] = { 1'b1, 8'h51, 8'h1f};
cfg[135] = { 1'b1, 8'h61, 8'h14};
cfg[136] = { 1'b1, 8'h71, 8'he};
cfg[137] = { 1'b1, 8'h81, 8'haf};
cfg[138] = { 1'b1, 8'h91, 8'h0};
cfg[139] = { 1'b1, 8'h39, 8'h1};
cfg[140] = { 1'b1, 8'h49, 8'h7f};
cfg[141] = { 1'b1, 8'h59, 8'h1f};
cfg[142] = { 1'b1, 8'h69, 8'h14};
cfg[143] = { 1'b1, 8'h79, 8'he};
cfg[144] = { 1'b1, 8'h89, 8'haf};
cfg[145] = { 1'b1, 8'h99, 8'h0};
cfg[146] = { 1'b1, 8'h35, 8'h1};
cfg[147] = { 1'b1, 8'h45, 8'h7f};
cfg[148] = { 1'b1, 8'h55, 8'h1f};
cfg[149] = { 1'b1, 8'h65, 8'h14};
cfg[150] = { 1'b1, 8'h75, 8'he};
cfg[151] = { 1'b1, 8'h85, 8'haf};
cfg[152] = { 1'b1, 8'h95, 8'h0};
cfg[153] = { 1'b1, 8'h3d, 8'h1};
cfg[154] = { 1'b1, 8'h4d, 8'h7f};
cfg[155] = { 1'b1, 8'h5d, 8'h1f};
cfg[156] = { 1'b1, 8'h6d, 8'h14};
cfg[157] = { 1'b1, 8'h7d, 8'he};
cfg[158] = { 1'b1, 8'h8d, 8'haf};
cfg[159] = { 1'b1, 8'h9d, 8'h0};
cfg[160] = { 1'b1, 8'ha2, 8'h0};
cfg[161] = { 1'b1, 8'ha6, 8'h24};
cfg[162] = { 1'b1, 8'hb2, 8'h7};
cfg[163] = { 1'b1, 8'hb6, 8'h0};
cfg[164] = { 1'b1, 8'h32, 8'h1};
cfg[165] = { 1'b1, 8'h42, 8'h7f};
cfg[166] = { 1'b1, 8'h52, 8'h1f};
cfg[167] = { 1'b1, 8'h62, 8'h14};
cfg[168] = { 1'b1, 8'h72, 8'he};
cfg[169] = { 1'b1, 8'h82, 8'haf};
cfg[170] = { 1'b1, 8'h92, 8'h0};
cfg[171] = { 1'b1, 8'h3a, 8'h1};
cfg[172] = { 1'b1, 8'h4a, 8'h7f};
cfg[173] = { 1'b1, 8'h5a, 8'h1f};
cfg[174] = { 1'b1, 8'h6a, 8'h14};
cfg[175] = { 1'b1, 8'h7a, 8'he};
cfg[176] = { 1'b1, 8'h8a, 8'haf};
cfg[177] = { 1'b1, 8'h9a, 8'h0};
cfg[178] = { 1'b1, 8'h36, 8'h1};
cfg[179] = { 1'b1, 8'h46, 8'h7f};
cfg[180] = { 1'b1, 8'h56, 8'h1f};
cfg[181] = { 1'b1, 8'h66, 8'h14};
cfg[182] = { 1'b1, 8'h76, 8'he};
cfg[183] = { 1'b1, 8'h86, 8'haf};
cfg[184] = { 1'b1, 8'h96, 8'h0};
cfg[185] = { 1'b1, 8'h3e, 8'h1};
cfg[186] = { 1'b1, 8'h4e, 8'h7f};
cfg[187] = { 1'b1, 8'h5e, 8'h1f};
cfg[188] = { 1'b1, 8'h6e, 8'h14};
cfg[189] = { 1'b1, 8'h7e, 8'he};
cfg[190] = { 1'b1, 8'h8e, 8'haf};
cfg[191] = { 1'b1, 8'h9e, 8'h0};
cfg[192] = { 1'b0, 8'h28, 8'hf0};
cfg[193] = { 1'b0, 8'h28, 8'hf1};
cfg[194] = { 1'b0, 8'h28, 8'hf2};
cfg[195] = { 1'b0, 8'h28, 8'hf4};
cfg[196] = { 1'b0, 8'h28, 8'hf5};
cfg[197] = { 1'b0, 8'h28, 8'hf6};
cfg[198] = { 1'b0, 8'h1, 8'hff};
cfg[199] = { 1'b0, 8'h28, 8'h0};
cfg[200] = { 1'b0, 8'h28, 8'h1};
cfg[201] = { 1'b0, 8'h28, 8'h2};
cfg[202] = { 1'b0, 8'h28, 8'h4};
cfg[203] = { 1'b0, 8'h28, 8'h5};
cfg[204] = { 1'b0, 8'h28, 8'h6};
cfg[205] = { 1'b0, 8'h1, 8'hff};
cfg[206] = { 1'b0, 8'hb0, 8'h7};
cfg[207] = { 1'b0, 8'hb0, 8'h27};
cfg[208] = { 1'b0, 8'hb1, 8'h7};
cfg[209] = { 1'b0, 8'hb1, 8'h27};
cfg[210] = { 1'b0, 8'hb2, 8'h7};
cfg[211] = { 1'b0, 8'hb2, 8'h27};
cfg[212] = { 1'b1, 8'hb0, 8'h7};
cfg[213] = { 1'b1, 8'hb0, 8'h27};
cfg[214] = { 1'b1, 8'hb1, 8'h7};
cfg[215] = { 1'b1, 8'hb1, 8'h27};
cfg[216] = { 1'b1, 8'hb2, 8'h7};
cfg[217] = { 1'b1, 8'hb2, 8'h27};
cfg[218] = { 1'b0, 8'h90, 8'h8};
cfg[219] = { 1'b0, 8'h40, 8'h0};
cfg[220] = { 1'b0, 8'h70, 8'h19};
cfg[221] = { 1'b0, 8'h60, 8'h1c};
cfg[222] = { 1'b0, 8'h98, 8'h9};
cfg[223] = { 1'b0, 8'h48, 8'h0};
cfg[224] = { 1'b0, 8'h78, 8'h19};
cfg[225] = { 1'b0, 8'h68, 8'h1c};
cfg[226] = { 1'b0, 8'h94, 8'ha};
cfg[227] = { 1'b0, 8'h44, 8'h0};
cfg[228] = { 1'b0, 8'h74, 8'h19};
cfg[229] = { 1'b0, 8'h64, 8'h1c};
cfg[230] = { 1'b0, 8'h9c, 8'hb};
cfg[231] = { 1'b0, 8'h4c, 8'h0};
cfg[232] = { 1'b0, 8'h7c, 8'h19};
cfg[233] = { 1'b0, 8'h6c, 8'h1c};
cfg[234] = { 1'b0, 8'h28, 8'hf0};
cfg[235] = { 1'b0, 8'h1, 8'hff};
cfg[236] = { 1'b0, 8'h1, 8'hff};
cfg[237] = { 1'b0, 8'h1, 8'hff};
cfg[238] = { 1'b0, 8'h1, 8'hff};
cfg[239] = { 1'b0, 8'h1, 8'hff};
cfg[240] = { 1'b0, 8'h1, 8'hff};
cfg[241] = { 1'b0, 8'h1, 8'hff};
cfg[242] = { 1'b0, 8'h28, 8'h0};
cfg[243] = { 1'b0, 8'h28, 8'h1};
cfg[244] = { 1'b0, 8'h28, 8'h2};
cfg[245] = { 1'b0, 8'h28, 8'h4};
cfg[246] = { 1'b0, 8'h28, 8'h5};
cfg[247] = { 1'b0, 8'h28, 8'h6};
cfg[248] = { 1'b0, 8'h91, 8'hc};
cfg[249] = { 1'b0, 8'h41, 8'h0};
cfg[250] = { 1'b0, 8'h71, 8'h19};
cfg[251] = { 1'b0, 8'h61, 8'h1c};
cfg[252] = { 1'b0, 8'h99, 8'hd};
cfg[253] = { 1'b0, 8'h49, 8'h0};
cfg[254] = { 1'b0, 8'h79, 8'h19};
cfg[255] = { 1'b0, 8'h69, 8'h1c};
cfg[256] = { 1'b0, 8'h95, 8'he};
cfg[257] = { 1'b0, 8'h45, 8'h0};
cfg[258] = { 1'b0, 8'h75, 8'h19};
cfg[259] = { 1'b0, 8'h65, 8'h1c};
cfg[260] = { 1'b0, 8'h9d, 8'hf};
cfg[261] = { 1'b0, 8'h4d, 8'h0};
cfg[262] = { 1'b0, 8'h7d, 8'h19};
cfg[263] = { 1'b0, 8'h6d, 8'h1c};
cfg[264] = { 1'b0, 8'h28, 8'hf1};
cfg[265] = { 1'b0, 8'h1, 8'hff};
cfg[266] = { 1'b0, 8'h1, 8'hff};
cfg[267] = { 1'b0, 8'h1, 8'hff};
cfg[268] = { 1'b0, 8'h1, 8'hff};
cfg[269] = { 1'b0, 8'h1, 8'hff};
cfg[270] = { 1'b0, 8'h1, 8'hff};
cfg[271] = { 1'b0, 8'h1, 8'hff};
cfg[272] = { 1'b0, 8'h28, 8'h0};
cfg[273] = { 1'b0, 8'h28, 8'h1};
cfg[274] = { 1'b0, 8'h28, 8'h2};
cfg[275] = { 1'b0, 8'h28, 8'h4};
cfg[276] = { 1'b0, 8'h28, 8'h5};
cfg[277] = { 1'b0, 8'h28, 8'h6};
cfg[278] = { 1'b0, 8'h92, 8'h8};
cfg[279] = { 1'b0, 8'h42, 8'h0};
cfg[280] = { 1'b0, 8'h72, 8'h19};
cfg[281] = { 1'b0, 8'h62, 8'h1c};
cfg[282] = { 1'b0, 8'h9a, 8'h9};
cfg[283] = { 1'b0, 8'h4a, 8'h0};
cfg[284] = { 1'b0, 8'h7a, 8'h19};
cfg[285] = { 1'b0, 8'h6a, 8'h1c};
cfg[286] = { 1'b0, 8'h96, 8'ha};
cfg[287] = { 1'b0, 8'h46, 8'h0};
cfg[288] = { 1'b0, 8'h76, 8'h19};
cfg[289] = { 1'b0, 8'h66, 8'h1c};
cfg[290] = { 1'b0, 8'h9e, 8'hb};
cfg[291] = { 1'b0, 8'h4e, 8'h0};
cfg[292] = { 1'b0, 8'h7e, 8'h19};
cfg[293] = { 1'b0, 8'h6e, 8'h1c};
cfg[294] = { 1'b0, 8'h28, 8'hf2};
cfg[295] = { 1'b0, 8'h1, 8'hff};
cfg[296] = { 1'b0, 8'h1, 8'hff};
cfg[297] = { 1'b0, 8'h1, 8'hff};
cfg[298] = { 1'b0, 8'h1, 8'hff};
cfg[299] = { 1'b0, 8'h1, 8'hff};
cfg[300] = { 1'b0, 8'h1, 8'hff};
cfg[301] = { 1'b0, 8'h1, 8'hff};
cfg[302] = { 1'b0, 8'h28, 8'h0};
cfg[303] = { 1'b0, 8'h28, 8'h1};
cfg[304] = { 1'b0, 8'h28, 8'h2};
cfg[305] = { 1'b0, 8'h28, 8'h4};
cfg[306] = { 1'b0, 8'h28, 8'h5};
cfg[307] = { 1'b0, 8'h28, 8'h6};
cfg[308] = { 1'b1, 8'h90, 8'hc};
cfg[309] = { 1'b1, 8'h40, 8'h0};
cfg[310] = { 1'b1, 8'h70, 8'h19};
cfg[311] = { 1'b1, 8'h60, 8'h1c};
cfg[312] = { 1'b1, 8'h98, 8'hd};
cfg[313] = { 1'b1, 8'h48, 8'h0};
cfg[314] = { 1'b1, 8'h78, 8'h19};
cfg[315] = { 1'b1, 8'h68, 8'h1c};
cfg[316] = { 1'b1, 8'h94, 8'he};
cfg[317] = { 1'b1, 8'h44, 8'h0};
cfg[318] = { 1'b1, 8'h74, 8'h19};
cfg[319] = { 1'b1, 8'h64, 8'h1c};
cfg[320] = { 1'b1, 8'h9c, 8'hf};
cfg[321] = { 1'b1, 8'h4c, 8'h0};
cfg[322] = { 1'b1, 8'h7c, 8'h19};
cfg[323] = { 1'b1, 8'h6c, 8'h1c};
cfg[324] = { 1'b0, 8'h28, 8'hf4};
cfg[325] = { 1'b0, 8'h1, 8'hff};
cfg[326] = { 1'b0, 8'h1, 8'hff};
cfg[327] = { 1'b0, 8'h1, 8'hff};
cfg[328] = { 1'b0, 8'h1, 8'hff};
cfg[329] = { 1'b0, 8'h1, 8'hff};
cfg[330] = { 1'b0, 8'h1, 8'hff};
cfg[331] = { 1'b0, 8'h1, 8'hff};
cfg[332] = { 1'b0, 8'h28, 8'h0};
cfg[333] = { 1'b0, 8'h28, 8'h1};
cfg[334] = { 1'b0, 8'h28, 8'h2};
cfg[335] = { 1'b0, 8'h28, 8'h4};
cfg[336] = { 1'b0, 8'h28, 8'h5};
cfg[337] = { 1'b0, 8'h28, 8'h6};
cfg[338] = { 1'b1, 8'h91, 8'h8};
cfg[339] = { 1'b1, 8'h41, 8'h0};
cfg[340] = { 1'b1, 8'h71, 8'h19};
cfg[341] = { 1'b1, 8'h61, 8'h1c};
cfg[342] = { 1'b1, 8'h99, 8'h9};
cfg[343] = { 1'b1, 8'h49, 8'h0};
cfg[344] = { 1'b1, 8'h79, 8'h19};
cfg[345] = { 1'b1, 8'h69, 8'h1c};
cfg[346] = { 1'b1, 8'h95, 8'ha};
cfg[347] = { 1'b1, 8'h45, 8'h0};
cfg[348] = { 1'b1, 8'h75, 8'h19};
cfg[349] = { 1'b1, 8'h65, 8'h1c};
cfg[350] = { 1'b1, 8'h9d, 8'hb};
cfg[351] = { 1'b1, 8'h4d, 8'h0};
cfg[352] = { 1'b1, 8'h7d, 8'h19};
cfg[353] = { 1'b1, 8'h6d, 8'h1c};
cfg[354] = { 1'b0, 8'h28, 8'hf5};
cfg[355] = { 1'b0, 8'h1, 8'hff};
cfg[356] = { 1'b0, 8'h1, 8'hff};
cfg[357] = { 1'b0, 8'h1, 8'hff};
cfg[358] = { 1'b0, 8'h1, 8'hff};
cfg[359] = { 1'b0, 8'h1, 8'hff};
cfg[360] = { 1'b0, 8'h1, 8'hff};
cfg[361] = { 1'b0, 8'h1, 8'hff};
cfg[362] = { 1'b0, 8'h28, 8'h0};
cfg[363] = { 1'b0, 8'h28, 8'h1};
cfg[364] = { 1'b0, 8'h28, 8'h2};
cfg[365] = { 1'b0, 8'h28, 8'h4};
cfg[366] = { 1'b0, 8'h28, 8'h5};
cfg[367] = { 1'b0, 8'h28, 8'h6};
cfg[368] = { 1'b1, 8'h92, 8'hc};
cfg[369] = { 1'b1, 8'h42, 8'h0};
cfg[370] = { 1'b1, 8'h72, 8'h19};
cfg[371] = { 1'b1, 8'h62, 8'h1c};
cfg[372] = { 1'b1, 8'h9a, 8'hd};
cfg[373] = { 1'b1, 8'h4a, 8'h0};
cfg[374] = { 1'b1, 8'h7a, 8'h19};
cfg[375] = { 1'b1, 8'h6a, 8'h1c};
cfg[376] = { 1'b1, 8'h96, 8'he};
cfg[377] = { 1'b1, 8'h46, 8'h0};
cfg[378] = { 1'b1, 8'h76, 8'h19};
cfg[379] = { 1'b1, 8'h66, 8'h1c};
cfg[380] = { 1'b1, 8'h9e, 8'hf};
cfg[381] = { 1'b1, 8'h4e, 8'h0};
cfg[382] = { 1'b1, 8'h7e, 8'h19};
cfg[383] = { 1'b1, 8'h6e, 8'h1c};
cfg[384] = { 1'b0, 8'h28, 8'hf6};
cfg[385] = { 1'b0, 8'h1, 8'hff};
cfg[386] = { 1'b0, 8'h1, 8'hff};
cfg[387] = { 1'b0, 8'h1, 8'hff};
cfg[388] = { 1'b0, 8'h1, 8'hff};
cfg[389] = { 1'b0, 8'h1, 8'hff};
cfg[390] = { 1'b0, 8'h1, 8'hff};
cfg[391] = { 1'b0, 8'h1, 8'hff};
cfg[392] = { 1'b0, 8'h28, 8'h0};
cfg[393] = { 1'b0, 8'h28, 8'h1};
cfg[394] = { 1'b0, 8'h28, 8'h2};
cfg[395] = { 1'b0, 8'h28, 8'h4};
cfg[396] = { 1'b0, 8'h28, 8'h5};
cfg[397] = { 1'b0, 8'h28, 8'h6};
cfg[398] = { 1'b0, 8'h90, 8'h0};
cfg[399] = { 1'b0, 8'h98, 8'h0};
cfg[400] = { 1'b0, 8'h94, 8'h0};
cfg[401] = { 1'b0, 8'h9c, 8'h0};
cfg[402] = { 1'b0, 8'h91, 8'h0};
cfg[403] = { 1'b0, 8'h99, 8'h0};
cfg[404] = { 1'b0, 8'h95, 8'h0};
cfg[405] = { 1'b0, 8'h9d, 8'h0};
cfg[406] = { 1'b0, 8'h92, 8'h0};
cfg[407] = { 1'b0, 8'h9a, 8'h0};
cfg[408] = { 1'b0, 8'h96, 8'h0};
cfg[409] = { 1'b0, 8'h9e, 8'h0};
cfg[410] = { 1'b1, 8'h90, 8'h0};
cfg[411] = { 1'b1, 8'h98, 8'h0};
cfg[412] = { 1'b1, 8'h94, 8'h0};
cfg[413] = { 1'b1, 8'h9c, 8'h0};
cfg[414] = { 1'b1, 8'h91, 8'h0};
cfg[415] = { 1'b1, 8'h99, 8'h0};
cfg[416] = { 1'b1, 8'h95, 8'h0};
cfg[417] = { 1'b1, 8'h9d, 8'h0};
cfg[418] = { 1'b1, 8'h92, 8'h0};
cfg[419] = { 1'b1, 8'h9a, 8'h0};
cfg[420] = { 1'b1, 8'h96, 8'h0};
cfg[421] = { 1'b1, 8'h9e, 8'h0};
cfg[422] = { 1'b0, 8'h40, 8'h0};
cfg[423] = { 1'b0, 8'h50, 8'h12};
cfg[424] = { 1'b0, 8'ha4, 8'hf};
cfg[425] = { 1'b0, 8'hb0, 8'h7};
cfg[426] = { 1'b0, 8'hb4, 8'hc0};
cfg[427] = { 1'b0, 8'h60, 8'h12};
cfg[428] = { 1'b0, 8'h70, 8'h12};
cfg[429] = { 1'b0, 8'h80, 8'h4f};
cfg[430] = { 1'b0, 8'h28, 8'h10};
cfg[431] = { 1'b0, 8'h1, 8'hff};
cfg[432] = { 1'b0, 8'h1, 8'hff};
cfg[433] = { 1'b0, 8'h1, 8'hff};
cfg[434] = { 1'b0, 8'h28, 8'h10};
cfg[435] = { 1'b0, 8'h1, 8'hff};
cfg[436] = { 1'b0, 8'h1, 8'hff};
cfg[437] = { 1'b0, 8'h1, 8'hff};
cfg[438] = { 1'b0, 8'h28, 8'h0};
cfg[439] = { 1'b0, 8'h1, 8'hff};
cfg[440] = { 1'b0, 8'h1, 8'hff};
cfg[441] = { 1'b0, 8'h1, 8'hff};
cfg[442] = { 1'b0, 8'h28, 8'h10};
cfg[443] = { 1'b0, 8'h1, 8'hff};
cfg[444] = { 1'b0, 8'h1, 8'hff};
cfg[445] = { 1'b0, 8'h1, 8'hff};
cfg[446] = { 1'b0, 8'h28, 8'h0};
cfg[447] = { 1'b0, 8'h1, 8'hff};
cfg[448] = { 1'b0, 8'h1, 8'hff};
cfg[449] = { 1'b0, 8'h1, 8'hff};
cfg[450] = { 1'b0, 8'h50, 8'h1f};
cfg[451] = { 1'b0, 8'h28, 8'h10};
cfg[452] = { 1'b0, 8'h1, 8'hff};
cfg[453] = { 1'b0, 8'h1, 8'hff};
cfg[454] = { 1'b0, 8'h1, 8'hff};
cfg[455] = { 1'b0, 8'h28, 8'h10};
cfg[456] = { 1'b0, 8'h1, 8'hff};
cfg[457] = { 1'b0, 8'h1, 8'hff};
cfg[458] = { 1'b0, 8'h1, 8'hff};
cfg[459] = { 1'b0, 8'h28, 8'h0};

cfg[460] = { 1'b0, 8'h0, 8'h00 }; // done
